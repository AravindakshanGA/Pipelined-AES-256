magic
tech sky130A
magscale 1 2
timestamp 1543373569
<< checkpaint >>
rect -1260 -1320 8139 26601
<< locali >>
rect 3988 25182 4004 25216
rect 4038 25182 4967 25216
rect 6284 25143 6861 25177
rect 4308 25070 4324 25104
rect 4358 25070 4857 25104
rect 4628 24980 4644 25014
rect 4678 24980 4967 25014
rect 4628 24756 4644 24790
rect 4678 24756 4967 24790
rect 4308 24666 4324 24700
rect 4358 24666 4857 24700
rect 6284 24593 6861 24627
rect 3908 24554 3924 24588
rect 3958 24554 4967 24588
rect 3828 24392 3844 24426
rect 3878 24392 4967 24426
rect 6284 24353 6861 24387
rect 4308 24280 4324 24314
rect 4358 24280 4857 24314
rect 4628 24190 4644 24224
rect 4678 24190 4967 24224
rect 4628 23966 4644 24000
rect 4678 23966 4967 24000
rect 4308 23876 4324 23910
rect 4358 23876 4857 23910
rect 6284 23803 6861 23837
rect 3748 23764 3764 23798
rect 3798 23764 4967 23798
rect 3988 23602 4004 23636
rect 4038 23602 4967 23636
rect 6284 23563 6861 23597
rect 4228 23490 4244 23524
rect 4278 23490 4857 23524
rect 4628 23400 4644 23434
rect 4678 23400 4967 23434
rect 4628 23176 4644 23210
rect 4678 23176 4967 23210
rect 4228 23086 4244 23120
rect 4278 23086 4857 23120
rect 6284 23013 6861 23047
rect 3908 22974 3924 23008
rect 3958 22974 4967 23008
rect 3828 22812 3844 22846
rect 3878 22812 4967 22846
rect 6284 22773 6861 22807
rect 4228 22700 4244 22734
rect 4278 22700 4857 22734
rect 4628 22610 4644 22644
rect 4678 22610 4967 22644
rect 4628 22386 4644 22420
rect 4678 22386 4967 22420
rect 4228 22296 4244 22330
rect 4278 22296 4857 22330
rect 6284 22223 6861 22257
rect 3748 22184 3764 22218
rect 3798 22184 4967 22218
rect 3988 22022 4004 22056
rect 4038 22022 4967 22056
rect 6284 21983 6861 22017
rect 4148 21910 4164 21944
rect 4198 21910 4857 21944
rect 4628 21820 4644 21854
rect 4678 21820 4967 21854
rect 4628 21596 4644 21630
rect 4678 21596 4967 21630
rect 4148 21506 4164 21540
rect 4198 21506 4857 21540
rect 6284 21433 6861 21467
rect 3908 21394 3924 21428
rect 3958 21394 4967 21428
rect 3828 21232 3844 21266
rect 3878 21232 4967 21266
rect 6284 21193 6861 21227
rect 4148 21120 4164 21154
rect 4198 21120 4857 21154
rect 4628 21030 4644 21064
rect 4678 21030 4967 21064
rect 4628 20806 4644 20840
rect 4678 20806 4967 20840
rect 4148 20716 4164 20750
rect 4198 20716 4857 20750
rect 6284 20643 6861 20677
rect 3748 20604 3764 20638
rect 3798 20604 4967 20638
rect 3988 20442 4004 20476
rect 4038 20442 4967 20476
rect 6284 20403 6861 20437
rect 4068 20330 4084 20364
rect 4118 20330 4857 20364
rect 4628 20240 4644 20274
rect 4678 20240 4967 20274
rect 4628 20016 4644 20050
rect 4678 20016 4967 20050
rect 4068 19926 4084 19960
rect 4118 19926 4857 19960
rect 6284 19853 6861 19887
rect 3908 19814 3924 19848
rect 3958 19814 4967 19848
rect 3828 19652 3844 19686
rect 3878 19652 4967 19686
rect 6284 19613 6861 19647
rect 4068 19540 4084 19574
rect 4118 19540 4857 19574
rect 4628 19450 4644 19484
rect 4678 19450 4967 19484
rect 4628 19226 4644 19260
rect 4678 19226 4967 19260
rect 4068 19136 4084 19170
rect 4118 19136 4857 19170
rect 6284 19063 6861 19097
rect 3748 19024 3764 19058
rect 3798 19024 4967 19058
rect 3988 18862 4004 18896
rect 4038 18862 4967 18896
rect 6284 18823 6861 18857
rect 4308 18750 4324 18784
rect 4358 18750 4857 18784
rect 4548 18660 4564 18694
rect 4598 18660 4967 18694
rect 4548 18436 4564 18470
rect 4598 18436 4967 18470
rect 4308 18346 4324 18380
rect 4358 18346 4857 18380
rect 6284 18273 6861 18307
rect 3908 18234 3924 18268
rect 3958 18234 4967 18268
rect 3828 18072 3844 18106
rect 3878 18072 4967 18106
rect 6284 18033 6861 18067
rect 4308 17960 4324 17994
rect 4358 17960 4857 17994
rect 4548 17870 4564 17904
rect 4598 17870 4967 17904
rect 4548 17646 4564 17680
rect 4598 17646 4967 17680
rect 4308 17556 4324 17590
rect 4358 17556 4857 17590
rect 6284 17483 6861 17517
rect 3748 17444 3764 17478
rect 3798 17444 4967 17478
rect 3988 17282 4004 17316
rect 4038 17282 4967 17316
rect 6284 17243 6861 17277
rect 4228 17170 4244 17204
rect 4278 17170 4857 17204
rect 4548 17080 4564 17114
rect 4598 17080 4967 17114
rect 4548 16856 4564 16890
rect 4598 16856 4967 16890
rect 4228 16766 4244 16800
rect 4278 16766 4857 16800
rect 6284 16693 6861 16727
rect 3908 16654 3924 16688
rect 3958 16654 4967 16688
rect 3828 16492 3844 16526
rect 3878 16492 4967 16526
rect 6284 16453 6861 16487
rect 4228 16380 4244 16414
rect 4278 16380 4857 16414
rect 4548 16290 4564 16324
rect 4598 16290 4967 16324
rect 4548 16066 4564 16100
rect 4598 16066 4967 16100
rect 4228 15976 4244 16010
rect 4278 15976 4857 16010
rect 6284 15903 6861 15937
rect 3748 15864 3764 15898
rect 3798 15864 4967 15898
rect 3988 15702 4004 15736
rect 4038 15702 4967 15736
rect 6284 15663 6861 15697
rect 4148 15590 4164 15624
rect 4198 15590 4857 15624
rect 4548 15500 4564 15534
rect 4598 15500 4967 15534
rect 4548 15276 4564 15310
rect 4598 15276 4967 15310
rect 4148 15186 4164 15220
rect 4198 15186 4857 15220
rect 6284 15113 6861 15147
rect 3908 15074 3924 15108
rect 3958 15074 4967 15108
rect 3828 14912 3844 14946
rect 3878 14912 4967 14946
rect 6284 14873 6861 14907
rect 4148 14800 4164 14834
rect 4198 14800 4857 14834
rect 4548 14710 4564 14744
rect 4598 14710 4967 14744
rect 4548 14486 4564 14520
rect 4598 14486 4967 14520
rect 4148 14396 4164 14430
rect 4198 14396 4857 14430
rect 6284 14323 6861 14357
rect 3748 14284 3764 14318
rect 3798 14284 4967 14318
rect 3988 14122 4004 14156
rect 4038 14122 4967 14156
rect 6284 14083 6861 14117
rect 4068 14010 4084 14044
rect 4118 14010 4857 14044
rect 4548 13920 4564 13954
rect 4598 13920 4967 13954
rect 4548 13696 4564 13730
rect 4598 13696 4967 13730
rect 4068 13606 4084 13640
rect 4118 13606 4857 13640
rect 6284 13533 6861 13567
rect 3908 13494 3924 13528
rect 3958 13494 4967 13528
rect 3828 13332 3844 13366
rect 3878 13332 4967 13366
rect 6284 13293 6861 13327
rect 4068 13220 4084 13254
rect 4118 13220 4857 13254
rect 4548 13130 4564 13164
rect 4598 13130 4967 13164
rect 4548 12906 4564 12940
rect 4598 12906 4967 12940
rect 4068 12816 4084 12850
rect 4118 12816 4857 12850
rect 6284 12743 6861 12777
rect 3748 12704 3764 12738
rect 3798 12704 4967 12738
rect 3988 12542 4004 12576
rect 4038 12542 4967 12576
rect 6284 12503 6861 12537
rect 4308 12430 4324 12464
rect 4358 12430 4857 12464
rect 4468 12340 4484 12374
rect 4518 12340 4967 12374
rect 4468 12116 4484 12150
rect 4518 12116 4967 12150
rect 4308 12026 4324 12060
rect 4358 12026 4857 12060
rect 6284 11953 6861 11987
rect 3908 11914 3924 11948
rect 3958 11914 4967 11948
rect 3828 11752 3844 11786
rect 3878 11752 4967 11786
rect 6284 11713 6861 11747
rect 4308 11640 4324 11674
rect 4358 11640 4857 11674
rect 4468 11550 4484 11584
rect 4518 11550 4967 11584
rect 4468 11326 4484 11360
rect 4518 11326 4967 11360
rect 4308 11236 4324 11270
rect 4358 11236 4857 11270
rect 6284 11163 6861 11197
rect 3748 11124 3764 11158
rect 3798 11124 4967 11158
rect 3988 10962 4004 10996
rect 4038 10962 4967 10996
rect 6284 10923 6861 10957
rect 4228 10850 4244 10884
rect 4278 10850 4857 10884
rect 4468 10760 4484 10794
rect 4518 10760 4967 10794
rect 4468 10536 4484 10570
rect 4518 10536 4967 10570
rect 4228 10446 4244 10480
rect 4278 10446 4857 10480
rect 6284 10373 6861 10407
rect 3908 10334 3924 10368
rect 3958 10334 4967 10368
rect 3828 10172 3844 10206
rect 3878 10172 4967 10206
rect 6284 10133 6861 10167
rect 4228 10060 4244 10094
rect 4278 10060 4857 10094
rect 4468 9970 4484 10004
rect 4518 9970 4967 10004
rect 4468 9746 4484 9780
rect 4518 9746 4967 9780
rect 4228 9656 4244 9690
rect 4278 9656 4857 9690
rect 6284 9583 6861 9617
rect 3748 9544 3764 9578
rect 3798 9544 4967 9578
rect 3988 9382 4004 9416
rect 4038 9382 4967 9416
rect 6284 9343 6861 9377
rect 4148 9270 4164 9304
rect 4198 9270 4857 9304
rect 4468 9180 4484 9214
rect 4518 9180 4967 9214
rect 4468 8956 4484 8990
rect 4518 8956 4967 8990
rect 4148 8866 4164 8900
rect 4198 8866 4857 8900
rect 6284 8793 6861 8827
rect 3908 8754 3924 8788
rect 3958 8754 4967 8788
rect 3828 8592 3844 8626
rect 3878 8592 4967 8626
rect 6284 8553 6861 8587
rect 4148 8480 4164 8514
rect 4198 8480 4857 8514
rect 4468 8390 4484 8424
rect 4518 8390 4967 8424
rect 4468 8166 4484 8200
rect 4518 8166 4967 8200
rect 4148 8076 4164 8110
rect 4198 8076 4857 8110
rect 6284 8003 6861 8037
rect 3748 7964 3764 7998
rect 3798 7964 4967 7998
rect 3988 7802 4004 7836
rect 4038 7802 4967 7836
rect 6284 7763 6861 7797
rect 4068 7690 4084 7724
rect 4118 7690 4857 7724
rect 4468 7600 4484 7634
rect 4518 7600 4967 7634
rect 4468 7376 4484 7410
rect 4518 7376 4967 7410
rect 4068 7286 4084 7320
rect 4118 7286 4857 7320
rect 6284 7213 6861 7247
rect 3908 7174 3924 7208
rect 3958 7174 4967 7208
rect 3828 7012 3844 7046
rect 3878 7012 4967 7046
rect 6284 6973 6861 7007
rect 4068 6900 4084 6934
rect 4118 6900 4857 6934
rect 4468 6810 4484 6844
rect 4518 6810 4967 6844
rect 4468 6586 4484 6620
rect 4518 6586 4967 6620
rect 4068 6496 4084 6530
rect 4118 6496 4857 6530
rect 6284 6423 6861 6457
rect 3748 6384 3764 6418
rect 3798 6384 4967 6418
rect 3670 6217 3704 6233
rect 3988 6222 4004 6256
rect 4038 6222 4967 6256
rect 6284 6183 6861 6217
rect 3670 6167 3704 6183
rect 4308 6110 4324 6144
rect 4358 6110 4857 6144
rect 4388 6020 4404 6054
rect 4438 6020 4967 6054
rect 4388 5796 4404 5830
rect 4438 5796 4967 5830
rect 4308 5706 4324 5740
rect 4358 5706 4857 5740
rect 3670 5667 3704 5683
rect 6284 5633 6861 5667
rect 3670 5617 3704 5633
rect 3908 5594 3924 5628
rect 3958 5594 4967 5628
rect 3670 5427 3704 5443
rect 3828 5432 3844 5466
rect 3878 5432 4967 5466
rect 6284 5393 6861 5427
rect 684 5377 718 5393
rect 3670 5377 3704 5393
rect 400 5343 416 5377
rect 450 5343 684 5377
rect 684 5327 718 5343
rect 4308 5320 4324 5354
rect 4358 5320 4857 5354
rect 4388 5230 4404 5264
rect 4438 5230 4967 5264
rect 4388 5006 4404 5040
rect 4438 5006 4967 5040
rect 604 4927 638 4943
rect 320 4893 336 4927
rect 370 4893 604 4927
rect 4308 4916 4324 4950
rect 4358 4916 4857 4950
rect 604 4877 638 4893
rect 3670 4877 3704 4893
rect 6284 4843 6861 4877
rect 3670 4827 3704 4843
rect 3748 4804 3764 4838
rect 3798 4804 4967 4838
rect 3988 4642 4004 4676
rect 4038 4642 4967 4676
rect 6284 4603 6861 4637
rect 4228 4530 4244 4564
rect 4278 4530 4857 4564
rect 4388 4440 4404 4474
rect 4438 4440 4967 4474
rect 4388 4216 4404 4250
rect 4438 4216 4967 4250
rect 4228 4126 4244 4160
rect 4278 4126 4857 4160
rect 6284 4053 6861 4087
rect 3908 4014 3924 4048
rect 3958 4014 4967 4048
rect 3670 3847 3704 3863
rect 3828 3852 3844 3886
rect 3878 3852 4967 3886
rect 6284 3813 6861 3847
rect 3670 3797 3704 3813
rect 4228 3740 4244 3774
rect 4278 3740 4857 3774
rect 4388 3650 4404 3684
rect 4438 3650 4967 3684
rect 4388 3426 4404 3460
rect 4438 3426 4967 3460
rect 4228 3336 4244 3370
rect 4278 3336 4857 3370
rect 3670 3297 3704 3313
rect 6284 3263 6861 3297
rect 3670 3247 3704 3263
rect 3748 3224 3764 3258
rect 3798 3224 4967 3258
rect 3670 3057 3704 3073
rect 3988 3062 4004 3096
rect 4038 3062 4967 3096
rect 6284 3023 6861 3057
rect 684 3007 718 3023
rect 3670 3007 3704 3023
rect 240 2973 256 3007
rect 290 2973 684 3007
rect 684 2957 718 2973
rect 4148 2950 4164 2984
rect 4198 2950 4857 2984
rect 4388 2860 4404 2894
rect 4438 2860 4967 2894
rect 4388 2636 4404 2670
rect 4438 2636 4967 2670
rect 604 2557 638 2573
rect 160 2523 176 2557
rect 210 2523 604 2557
rect 4148 2546 4164 2580
rect 4198 2546 4857 2580
rect 604 2507 638 2523
rect 3670 2507 3704 2523
rect 6284 2473 6861 2507
rect 3670 2457 3704 2473
rect 3908 2434 3924 2468
rect 3958 2434 4967 2468
rect 3828 2272 3844 2306
rect 3878 2272 4967 2306
rect 6284 2233 6861 2267
rect 4148 2160 4164 2194
rect 4198 2160 4857 2194
rect 4388 2070 4404 2104
rect 4438 2070 4967 2104
rect 4388 1846 4404 1880
rect 4438 1846 4967 1880
rect 4148 1756 4164 1790
rect 4198 1756 4857 1790
rect 6284 1683 6861 1717
rect 3748 1644 3764 1678
rect 3798 1644 4967 1678
rect 3670 1477 3704 1493
rect 3988 1482 4004 1516
rect 4038 1482 4967 1516
rect 6284 1443 6861 1477
rect 3670 1427 3704 1443
rect 4068 1370 4084 1404
rect 4118 1370 4857 1404
rect 4388 1280 4404 1314
rect 4438 1280 4967 1314
rect 4388 1056 4404 1090
rect 4438 1056 4967 1090
rect 4068 966 4084 1000
rect 4118 966 4857 1000
rect 3670 927 3704 943
rect 6284 893 6861 927
rect 3670 877 3704 893
rect 3908 854 3924 888
rect 3958 854 4967 888
rect 3670 687 3704 703
rect 3828 692 3844 726
rect 3878 692 4967 726
rect 6284 653 6861 687
rect 684 637 718 653
rect 3670 637 3704 653
rect 80 603 96 637
rect 130 603 684 637
rect 684 587 718 603
rect 4068 580 4084 614
rect 4118 580 4857 614
rect 4388 490 4404 524
rect 4438 490 4967 524
rect 4388 266 4404 300
rect 4438 266 4967 300
rect 604 187 638 203
rect 0 153 16 187
rect 50 153 604 187
rect 4068 176 4084 210
rect 4118 176 4857 210
rect 604 137 638 153
rect 3670 137 3704 153
rect 6284 103 6861 137
rect 3670 87 3704 103
rect 3748 64 3764 98
rect 3798 64 4967 98
<< viali >>
rect 4004 25182 4038 25216
rect 4324 25070 4358 25104
rect 4644 24980 4678 25014
rect 4644 24756 4678 24790
rect 4324 24666 4358 24700
rect 3924 24554 3958 24588
rect 3844 24392 3878 24426
rect 4324 24280 4358 24314
rect 4644 24190 4678 24224
rect 4644 23966 4678 24000
rect 4324 23876 4358 23910
rect 3764 23764 3798 23798
rect 4004 23602 4038 23636
rect 4244 23490 4278 23524
rect 4644 23400 4678 23434
rect 4644 23176 4678 23210
rect 4244 23086 4278 23120
rect 3924 22974 3958 23008
rect 3844 22812 3878 22846
rect 4244 22700 4278 22734
rect 4644 22610 4678 22644
rect 4644 22386 4678 22420
rect 4244 22296 4278 22330
rect 3764 22184 3798 22218
rect 4004 22022 4038 22056
rect 4164 21910 4198 21944
rect 4644 21820 4678 21854
rect 4644 21596 4678 21630
rect 4164 21506 4198 21540
rect 3924 21394 3958 21428
rect 3844 21232 3878 21266
rect 4164 21120 4198 21154
rect 4644 21030 4678 21064
rect 4644 20806 4678 20840
rect 4164 20716 4198 20750
rect 3764 20604 3798 20638
rect 4004 20442 4038 20476
rect 4084 20330 4118 20364
rect 4644 20240 4678 20274
rect 4644 20016 4678 20050
rect 4084 19926 4118 19960
rect 3924 19814 3958 19848
rect 3844 19652 3878 19686
rect 4084 19540 4118 19574
rect 4644 19450 4678 19484
rect 4644 19226 4678 19260
rect 4084 19136 4118 19170
rect 3764 19024 3798 19058
rect 4004 18862 4038 18896
rect 4324 18750 4358 18784
rect 4564 18660 4598 18694
rect 4564 18436 4598 18470
rect 4324 18346 4358 18380
rect 3924 18234 3958 18268
rect 3844 18072 3878 18106
rect 4324 17960 4358 17994
rect 4564 17870 4598 17904
rect 4564 17646 4598 17680
rect 4324 17556 4358 17590
rect 3764 17444 3798 17478
rect 4004 17282 4038 17316
rect 4244 17170 4278 17204
rect 4564 17080 4598 17114
rect 4564 16856 4598 16890
rect 4244 16766 4278 16800
rect 3924 16654 3958 16688
rect 3844 16492 3878 16526
rect 4244 16380 4278 16414
rect 4564 16290 4598 16324
rect 4564 16066 4598 16100
rect 4244 15976 4278 16010
rect 3764 15864 3798 15898
rect 4004 15702 4038 15736
rect 4164 15590 4198 15624
rect 4564 15500 4598 15534
rect 4564 15276 4598 15310
rect 4164 15186 4198 15220
rect 3924 15074 3958 15108
rect 3844 14912 3878 14946
rect 4164 14800 4198 14834
rect 4564 14710 4598 14744
rect 4564 14486 4598 14520
rect 4164 14396 4198 14430
rect 3764 14284 3798 14318
rect 4004 14122 4038 14156
rect 4084 14010 4118 14044
rect 4564 13920 4598 13954
rect 4564 13696 4598 13730
rect 4084 13606 4118 13640
rect 3924 13494 3958 13528
rect 3844 13332 3878 13366
rect 4084 13220 4118 13254
rect 4564 13130 4598 13164
rect 4564 12906 4598 12940
rect 4084 12816 4118 12850
rect 3764 12704 3798 12738
rect 4004 12542 4038 12576
rect 4324 12430 4358 12464
rect 4484 12340 4518 12374
rect 4484 12116 4518 12150
rect 4324 12026 4358 12060
rect 3924 11914 3958 11948
rect 3844 11752 3878 11786
rect 4324 11640 4358 11674
rect 4484 11550 4518 11584
rect 4484 11326 4518 11360
rect 4324 11236 4358 11270
rect 3764 11124 3798 11158
rect 4004 10962 4038 10996
rect 4244 10850 4278 10884
rect 4484 10760 4518 10794
rect 4484 10536 4518 10570
rect 4244 10446 4278 10480
rect 3924 10334 3958 10368
rect 3844 10172 3878 10206
rect 4244 10060 4278 10094
rect 4484 9970 4518 10004
rect 4484 9746 4518 9780
rect 4244 9656 4278 9690
rect 3764 9544 3798 9578
rect 4004 9382 4038 9416
rect 4164 9270 4198 9304
rect 4484 9180 4518 9214
rect 4484 8956 4518 8990
rect 4164 8866 4198 8900
rect 3924 8754 3958 8788
rect 3844 8592 3878 8626
rect 4164 8480 4198 8514
rect 4484 8390 4518 8424
rect 4484 8166 4518 8200
rect 4164 8076 4198 8110
rect 3764 7964 3798 7998
rect 4004 7802 4038 7836
rect 4084 7690 4118 7724
rect 4484 7600 4518 7634
rect 4484 7376 4518 7410
rect 4084 7286 4118 7320
rect 3924 7174 3958 7208
rect 3844 7012 3878 7046
rect 4084 6900 4118 6934
rect 4484 6810 4518 6844
rect 4484 6586 4518 6620
rect 4084 6496 4118 6530
rect 3764 6384 3798 6418
rect 4004 6222 4038 6256
rect 3670 6183 3704 6217
rect 4324 6110 4358 6144
rect 4404 6020 4438 6054
rect 4404 5796 4438 5830
rect 4324 5706 4358 5740
rect 3670 5633 3704 5667
rect 3924 5594 3958 5628
rect 3844 5432 3878 5466
rect 3670 5393 3704 5427
rect 416 5343 450 5377
rect 684 5343 718 5377
rect 4324 5320 4358 5354
rect 4404 5230 4438 5264
rect 4404 5006 4438 5040
rect 336 4893 370 4927
rect 604 4893 638 4927
rect 4324 4916 4358 4950
rect 3670 4843 3704 4877
rect 3764 4804 3798 4838
rect 4004 4642 4038 4676
rect 4244 4530 4278 4564
rect 4404 4440 4438 4474
rect 4404 4216 4438 4250
rect 4244 4126 4278 4160
rect 3924 4014 3958 4048
rect 3844 3852 3878 3886
rect 3670 3813 3704 3847
rect 4244 3740 4278 3774
rect 4404 3650 4438 3684
rect 4404 3426 4438 3460
rect 4244 3336 4278 3370
rect 3670 3263 3704 3297
rect 3764 3224 3798 3258
rect 4004 3062 4038 3096
rect 3670 3023 3704 3057
rect 256 2973 290 3007
rect 684 2973 718 3007
rect 4164 2950 4198 2984
rect 4404 2860 4438 2894
rect 4404 2636 4438 2670
rect 176 2523 210 2557
rect 604 2523 638 2557
rect 4164 2546 4198 2580
rect 3670 2473 3704 2507
rect 3924 2434 3958 2468
rect 3844 2272 3878 2306
rect 4164 2160 4198 2194
rect 4404 2070 4438 2104
rect 4404 1846 4438 1880
rect 4164 1756 4198 1790
rect 3764 1644 3798 1678
rect 4004 1482 4038 1516
rect 3670 1443 3704 1477
rect 4084 1370 4118 1404
rect 4404 1280 4438 1314
rect 4404 1056 4438 1090
rect 4084 966 4118 1000
rect 3670 893 3704 927
rect 3924 854 3958 888
rect 3844 692 3878 726
rect 3670 653 3704 687
rect 96 603 130 637
rect 684 603 718 637
rect 4084 580 4118 614
rect 4404 490 4438 524
rect 4404 266 4438 300
rect 16 153 50 187
rect 604 153 638 187
rect 4084 176 4118 210
rect 3670 103 3704 137
rect 3764 64 3798 98
<< metal1 >>
rect 3767 23810 3795 25308
rect 3847 24438 3875 25308
rect 3927 24600 3955 25308
rect 4007 25228 4035 25308
rect 3998 25216 4044 25228
rect 3998 25182 4004 25216
rect 4038 25182 4044 25216
rect 3998 25170 4044 25182
rect 3918 24588 3964 24600
rect 3918 24554 3924 24588
rect 3958 24554 3964 24588
rect 3918 24542 3964 24554
rect 3838 24426 3884 24438
rect 3838 24392 3844 24426
rect 3878 24392 3884 24426
rect 3838 24380 3884 24392
rect 3758 23798 3804 23810
rect 3758 23764 3764 23798
rect 3798 23764 3804 23798
rect 3758 23752 3804 23764
rect 3767 22230 3795 23752
rect 3847 22858 3875 24380
rect 3927 23020 3955 24542
rect 4007 23648 4035 25170
rect 3998 23636 4044 23648
rect 3998 23602 4004 23636
rect 4038 23602 4044 23636
rect 3998 23590 4044 23602
rect 3918 23008 3964 23020
rect 3918 22974 3924 23008
rect 3958 22974 3964 23008
rect 3918 22962 3964 22974
rect 3838 22846 3884 22858
rect 3838 22812 3844 22846
rect 3878 22812 3884 22846
rect 3838 22800 3884 22812
rect 3758 22218 3804 22230
rect 3758 22184 3764 22218
rect 3798 22184 3804 22218
rect 3758 22172 3804 22184
rect 3767 20650 3795 22172
rect 3847 21278 3875 22800
rect 3927 21440 3955 22962
rect 4007 22068 4035 23590
rect 3998 22056 4044 22068
rect 3998 22022 4004 22056
rect 4038 22022 4044 22056
rect 3998 22010 4044 22022
rect 3918 21428 3964 21440
rect 3918 21394 3924 21428
rect 3958 21394 3964 21428
rect 3918 21382 3964 21394
rect 3838 21266 3884 21278
rect 3838 21232 3844 21266
rect 3878 21232 3884 21266
rect 3838 21220 3884 21232
rect 3758 20638 3804 20650
rect 3758 20604 3764 20638
rect 3798 20604 3804 20638
rect 3758 20592 3804 20604
rect 3767 19070 3795 20592
rect 3847 19698 3875 21220
rect 3927 19860 3955 21382
rect 4007 20488 4035 22010
rect 3998 20476 4044 20488
rect 3998 20442 4004 20476
rect 4038 20442 4044 20476
rect 3998 20430 4044 20442
rect 3918 19848 3964 19860
rect 3918 19814 3924 19848
rect 3958 19814 3964 19848
rect 3918 19802 3964 19814
rect 3838 19686 3884 19698
rect 3838 19652 3844 19686
rect 3878 19652 3884 19686
rect 3838 19640 3884 19652
rect 3758 19058 3804 19070
rect 3758 19024 3764 19058
rect 3798 19024 3804 19058
rect 3758 19012 3804 19024
rect 3767 17490 3795 19012
rect 3847 18118 3875 19640
rect 3927 18280 3955 19802
rect 4007 18908 4035 20430
rect 4087 20376 4115 25308
rect 4167 21956 4195 25308
rect 4247 23536 4275 25308
rect 4327 25116 4355 25308
rect 4318 25104 4364 25116
rect 4318 25070 4324 25104
rect 4358 25070 4364 25104
rect 4318 25058 4364 25070
rect 4327 24712 4355 25058
rect 4318 24700 4364 24712
rect 4318 24666 4324 24700
rect 4358 24666 4364 24700
rect 4318 24654 4364 24666
rect 4327 24326 4355 24654
rect 4318 24314 4364 24326
rect 4318 24280 4324 24314
rect 4358 24280 4364 24314
rect 4318 24268 4364 24280
rect 4327 23922 4355 24268
rect 4318 23910 4364 23922
rect 4318 23876 4324 23910
rect 4358 23876 4364 23910
rect 4318 23864 4364 23876
rect 4238 23524 4284 23536
rect 4238 23490 4244 23524
rect 4278 23490 4284 23524
rect 4238 23478 4284 23490
rect 4247 23132 4275 23478
rect 4238 23120 4284 23132
rect 4238 23086 4244 23120
rect 4278 23086 4284 23120
rect 4238 23074 4284 23086
rect 4247 22746 4275 23074
rect 4238 22734 4284 22746
rect 4238 22700 4244 22734
rect 4278 22700 4284 22734
rect 4238 22688 4284 22700
rect 4247 22342 4275 22688
rect 4238 22330 4284 22342
rect 4238 22296 4244 22330
rect 4278 22296 4284 22330
rect 4238 22284 4284 22296
rect 4158 21944 4204 21956
rect 4158 21910 4164 21944
rect 4198 21910 4204 21944
rect 4158 21898 4204 21910
rect 4167 21552 4195 21898
rect 4158 21540 4204 21552
rect 4158 21506 4164 21540
rect 4198 21506 4204 21540
rect 4158 21494 4204 21506
rect 4167 21166 4195 21494
rect 4158 21154 4204 21166
rect 4158 21120 4164 21154
rect 4198 21120 4204 21154
rect 4158 21108 4204 21120
rect 4167 20762 4195 21108
rect 4158 20750 4204 20762
rect 4158 20716 4164 20750
rect 4198 20716 4204 20750
rect 4158 20704 4204 20716
rect 4078 20364 4124 20376
rect 4078 20330 4084 20364
rect 4118 20330 4124 20364
rect 4078 20318 4124 20330
rect 4087 19972 4115 20318
rect 4078 19960 4124 19972
rect 4078 19926 4084 19960
rect 4118 19926 4124 19960
rect 4078 19914 4124 19926
rect 4087 19586 4115 19914
rect 4078 19574 4124 19586
rect 4078 19540 4084 19574
rect 4118 19540 4124 19574
rect 4078 19528 4124 19540
rect 4087 19182 4115 19528
rect 4078 19170 4124 19182
rect 4078 19136 4084 19170
rect 4118 19136 4124 19170
rect 4078 19124 4124 19136
rect 3998 18896 4044 18908
rect 3998 18862 4004 18896
rect 4038 18862 4044 18896
rect 3998 18850 4044 18862
rect 3918 18268 3964 18280
rect 3918 18234 3924 18268
rect 3958 18234 3964 18268
rect 3918 18222 3964 18234
rect 3838 18106 3884 18118
rect 3838 18072 3844 18106
rect 3878 18072 3884 18106
rect 3838 18060 3884 18072
rect 3758 17478 3804 17490
rect 3758 17444 3764 17478
rect 3798 17444 3804 17478
rect 3758 17432 3804 17444
rect 3767 15910 3795 17432
rect 3847 16538 3875 18060
rect 3927 16700 3955 18222
rect 4007 17328 4035 18850
rect 3998 17316 4044 17328
rect 3998 17282 4004 17316
rect 4038 17282 4044 17316
rect 3998 17270 4044 17282
rect 3918 16688 3964 16700
rect 3918 16654 3924 16688
rect 3958 16654 3964 16688
rect 3918 16642 3964 16654
rect 3838 16526 3884 16538
rect 3838 16492 3844 16526
rect 3878 16492 3884 16526
rect 3838 16480 3884 16492
rect 3758 15898 3804 15910
rect 3758 15864 3764 15898
rect 3798 15864 3804 15898
rect 3758 15852 3804 15864
rect 3767 14330 3795 15852
rect 3847 14958 3875 16480
rect 3927 15120 3955 16642
rect 4007 15748 4035 17270
rect 3998 15736 4044 15748
rect 3998 15702 4004 15736
rect 4038 15702 4044 15736
rect 3998 15690 4044 15702
rect 3918 15108 3964 15120
rect 3918 15074 3924 15108
rect 3958 15074 3964 15108
rect 3918 15062 3964 15074
rect 3838 14946 3884 14958
rect 3838 14912 3844 14946
rect 3878 14912 3884 14946
rect 3838 14900 3884 14912
rect 3758 14318 3804 14330
rect 3758 14284 3764 14318
rect 3798 14284 3804 14318
rect 3758 14272 3804 14284
rect 3767 12750 3795 14272
rect 3847 13378 3875 14900
rect 3927 13540 3955 15062
rect 4007 14168 4035 15690
rect 3998 14156 4044 14168
rect 3998 14122 4004 14156
rect 4038 14122 4044 14156
rect 3998 14110 4044 14122
rect 3918 13528 3964 13540
rect 3918 13494 3924 13528
rect 3958 13494 3964 13528
rect 3918 13482 3964 13494
rect 3838 13366 3884 13378
rect 3838 13332 3844 13366
rect 3878 13332 3884 13366
rect 3838 13320 3884 13332
rect 3758 12738 3804 12750
rect 3758 12704 3764 12738
rect 3798 12704 3804 12738
rect 3758 12692 3804 12704
rect 3767 11170 3795 12692
rect 3847 11798 3875 13320
rect 3927 11960 3955 13482
rect 4007 12588 4035 14110
rect 4087 14056 4115 19124
rect 4167 15636 4195 20704
rect 4247 17216 4275 22284
rect 4327 18796 4355 23864
rect 4318 18784 4364 18796
rect 4318 18750 4324 18784
rect 4358 18750 4364 18784
rect 4318 18738 4364 18750
rect 4327 18392 4355 18738
rect 4318 18380 4364 18392
rect 4318 18346 4324 18380
rect 4358 18346 4364 18380
rect 4318 18334 4364 18346
rect 4327 18006 4355 18334
rect 4318 17994 4364 18006
rect 4318 17960 4324 17994
rect 4358 17960 4364 17994
rect 4318 17948 4364 17960
rect 4327 17602 4355 17948
rect 4318 17590 4364 17602
rect 4318 17556 4324 17590
rect 4358 17556 4364 17590
rect 4318 17544 4364 17556
rect 4238 17204 4284 17216
rect 4238 17170 4244 17204
rect 4278 17170 4284 17204
rect 4238 17158 4284 17170
rect 4247 16812 4275 17158
rect 4238 16800 4284 16812
rect 4238 16766 4244 16800
rect 4278 16766 4284 16800
rect 4238 16754 4284 16766
rect 4247 16426 4275 16754
rect 4238 16414 4284 16426
rect 4238 16380 4244 16414
rect 4278 16380 4284 16414
rect 4238 16368 4284 16380
rect 4247 16022 4275 16368
rect 4238 16010 4284 16022
rect 4238 15976 4244 16010
rect 4278 15976 4284 16010
rect 4238 15964 4284 15976
rect 4158 15624 4204 15636
rect 4158 15590 4164 15624
rect 4198 15590 4204 15624
rect 4158 15578 4204 15590
rect 4167 15232 4195 15578
rect 4158 15220 4204 15232
rect 4158 15186 4164 15220
rect 4198 15186 4204 15220
rect 4158 15174 4204 15186
rect 4167 14846 4195 15174
rect 4158 14834 4204 14846
rect 4158 14800 4164 14834
rect 4198 14800 4204 14834
rect 4158 14788 4204 14800
rect 4167 14442 4195 14788
rect 4158 14430 4204 14442
rect 4158 14396 4164 14430
rect 4198 14396 4204 14430
rect 4158 14384 4204 14396
rect 4078 14044 4124 14056
rect 4078 14010 4084 14044
rect 4118 14010 4124 14044
rect 4078 13998 4124 14010
rect 4087 13652 4115 13998
rect 4078 13640 4124 13652
rect 4078 13606 4084 13640
rect 4118 13606 4124 13640
rect 4078 13594 4124 13606
rect 4087 13266 4115 13594
rect 4078 13254 4124 13266
rect 4078 13220 4084 13254
rect 4118 13220 4124 13254
rect 4078 13208 4124 13220
rect 4087 12862 4115 13208
rect 4078 12850 4124 12862
rect 4078 12816 4084 12850
rect 4118 12816 4124 12850
rect 4078 12804 4124 12816
rect 3998 12576 4044 12588
rect 3998 12542 4004 12576
rect 4038 12542 4044 12576
rect 3998 12530 4044 12542
rect 3918 11948 3964 11960
rect 3918 11914 3924 11948
rect 3958 11914 3964 11948
rect 3918 11902 3964 11914
rect 3838 11786 3884 11798
rect 3838 11752 3844 11786
rect 3878 11752 3884 11786
rect 3838 11740 3884 11752
rect 3758 11158 3804 11170
rect 3758 11124 3764 11158
rect 3798 11124 3804 11158
rect 3758 11112 3804 11124
rect 3767 9590 3795 11112
rect 3847 10218 3875 11740
rect 3927 10380 3955 11902
rect 4007 11008 4035 12530
rect 3998 10996 4044 11008
rect 3998 10962 4004 10996
rect 4038 10962 4044 10996
rect 3998 10950 4044 10962
rect 3918 10368 3964 10380
rect 3918 10334 3924 10368
rect 3958 10334 3964 10368
rect 3918 10322 3964 10334
rect 3838 10206 3884 10218
rect 3838 10172 3844 10206
rect 3878 10172 3884 10206
rect 3838 10160 3884 10172
rect 3758 9578 3804 9590
rect 3758 9544 3764 9578
rect 3798 9544 3804 9578
rect 3758 9532 3804 9544
rect 3767 8010 3795 9532
rect 3847 8638 3875 10160
rect 3927 8800 3955 10322
rect 4007 9428 4035 10950
rect 3998 9416 4044 9428
rect 3998 9382 4004 9416
rect 4038 9382 4044 9416
rect 3998 9370 4044 9382
rect 3918 8788 3964 8800
rect 3918 8754 3924 8788
rect 3958 8754 3964 8788
rect 3918 8742 3964 8754
rect 3838 8626 3884 8638
rect 3838 8592 3844 8626
rect 3878 8592 3884 8626
rect 3838 8580 3884 8592
rect 3758 7998 3804 8010
rect 3758 7964 3764 7998
rect 3798 7964 3804 7998
rect 3758 7952 3804 7964
rect 3767 6430 3795 7952
rect 3847 7058 3875 8580
rect 3927 7220 3955 8742
rect 4007 7848 4035 9370
rect 3998 7836 4044 7848
rect 3998 7802 4004 7836
rect 4038 7802 4044 7836
rect 3998 7790 4044 7802
rect 3918 7208 3964 7220
rect 3918 7174 3924 7208
rect 3958 7174 3964 7208
rect 3918 7162 3964 7174
rect 3838 7046 3884 7058
rect 3838 7012 3844 7046
rect 3878 7012 3884 7046
rect 3838 7000 3884 7012
rect 3758 6418 3804 6430
rect 3758 6384 3764 6418
rect 3798 6384 3804 6418
rect 3758 6372 3804 6384
rect 19 199 47 6320
rect 99 649 127 6320
rect 179 2569 207 6320
rect 259 3019 287 6320
rect 339 4939 367 6320
rect 419 5389 447 6320
rect 3655 6174 3661 6226
rect 3713 6174 3719 6226
rect 3655 5624 3661 5676
rect 3713 5624 3719 5676
rect 410 5377 456 5389
rect 3655 5384 3661 5436
rect 3713 5384 3719 5436
rect 410 5343 416 5377
rect 450 5343 456 5377
rect 410 5331 456 5343
rect 672 5377 730 5383
rect 672 5343 684 5377
rect 718 5343 730 5377
rect 672 5337 730 5343
rect 330 4927 376 4939
rect 330 4893 336 4927
rect 370 4893 376 4927
rect 330 4881 376 4893
rect 250 3007 296 3019
rect 250 2973 256 3007
rect 290 2973 296 3007
rect 250 2961 296 2973
rect 170 2557 216 2569
rect 170 2523 176 2557
rect 210 2523 216 2557
rect 170 2511 216 2523
rect 90 637 136 649
rect 90 603 96 637
rect 130 603 136 637
rect 90 591 136 603
rect 10 187 56 199
rect 10 153 16 187
rect 50 153 56 187
rect 10 141 56 153
rect 19 0 47 141
rect 99 0 127 591
rect 179 0 207 2511
rect 259 0 287 2961
rect 339 0 367 4881
rect 419 0 447 5331
rect 592 4927 650 4933
rect 592 4893 604 4927
rect 638 4893 650 4927
rect 592 4887 650 4893
rect 3655 4834 3661 4886
rect 3713 4834 3719 4886
rect 3767 4850 3795 6372
rect 3847 5478 3875 7000
rect 3927 5640 3955 7162
rect 4007 6268 4035 7790
rect 4087 7736 4115 12804
rect 4167 9316 4195 14384
rect 4247 10896 4275 15964
rect 4327 12476 4355 17544
rect 4318 12464 4364 12476
rect 4318 12430 4324 12464
rect 4358 12430 4364 12464
rect 4318 12418 4364 12430
rect 4327 12072 4355 12418
rect 4318 12060 4364 12072
rect 4318 12026 4324 12060
rect 4358 12026 4364 12060
rect 4318 12014 4364 12026
rect 4327 11686 4355 12014
rect 4318 11674 4364 11686
rect 4318 11640 4324 11674
rect 4358 11640 4364 11674
rect 4318 11628 4364 11640
rect 4327 11282 4355 11628
rect 4318 11270 4364 11282
rect 4318 11236 4324 11270
rect 4358 11236 4364 11270
rect 4318 11224 4364 11236
rect 4238 10884 4284 10896
rect 4238 10850 4244 10884
rect 4278 10850 4284 10884
rect 4238 10838 4284 10850
rect 4247 10492 4275 10838
rect 4238 10480 4284 10492
rect 4238 10446 4244 10480
rect 4278 10446 4284 10480
rect 4238 10434 4284 10446
rect 4247 10106 4275 10434
rect 4238 10094 4284 10106
rect 4238 10060 4244 10094
rect 4278 10060 4284 10094
rect 4238 10048 4284 10060
rect 4247 9702 4275 10048
rect 4238 9690 4284 9702
rect 4238 9656 4244 9690
rect 4278 9656 4284 9690
rect 4238 9644 4284 9656
rect 4158 9304 4204 9316
rect 4158 9270 4164 9304
rect 4198 9270 4204 9304
rect 4158 9258 4204 9270
rect 4167 8912 4195 9258
rect 4158 8900 4204 8912
rect 4158 8866 4164 8900
rect 4198 8866 4204 8900
rect 4158 8854 4204 8866
rect 4167 8526 4195 8854
rect 4158 8514 4204 8526
rect 4158 8480 4164 8514
rect 4198 8480 4204 8514
rect 4158 8468 4204 8480
rect 4167 8122 4195 8468
rect 4158 8110 4204 8122
rect 4158 8076 4164 8110
rect 4198 8076 4204 8110
rect 4158 8064 4204 8076
rect 4078 7724 4124 7736
rect 4078 7690 4084 7724
rect 4118 7690 4124 7724
rect 4078 7678 4124 7690
rect 4087 7332 4115 7678
rect 4078 7320 4124 7332
rect 4078 7286 4084 7320
rect 4118 7286 4124 7320
rect 4078 7274 4124 7286
rect 4087 6946 4115 7274
rect 4078 6934 4124 6946
rect 4078 6900 4084 6934
rect 4118 6900 4124 6934
rect 4078 6888 4124 6900
rect 4087 6542 4115 6888
rect 4078 6530 4124 6542
rect 4078 6496 4084 6530
rect 4118 6496 4124 6530
rect 4078 6484 4124 6496
rect 3998 6256 4044 6268
rect 3998 6222 4004 6256
rect 4038 6222 4044 6256
rect 3998 6210 4044 6222
rect 3918 5628 3964 5640
rect 3918 5594 3924 5628
rect 3958 5594 3964 5628
rect 3918 5582 3964 5594
rect 3838 5466 3884 5478
rect 3838 5432 3844 5466
rect 3878 5432 3884 5466
rect 3838 5420 3884 5432
rect 3758 4838 3804 4850
rect 3758 4804 3764 4838
rect 3798 4804 3804 4838
rect 3758 4792 3804 4804
rect 3655 3804 3661 3856
rect 3713 3804 3719 3856
rect 3655 3254 3661 3306
rect 3713 3254 3719 3306
rect 3767 3270 3795 4792
rect 3847 3898 3875 5420
rect 3927 4060 3955 5582
rect 4007 4688 4035 6210
rect 3998 4676 4044 4688
rect 3998 4642 4004 4676
rect 4038 4642 4044 4676
rect 3998 4630 4044 4642
rect 3918 4048 3964 4060
rect 3918 4014 3924 4048
rect 3958 4014 3964 4048
rect 3918 4002 3964 4014
rect 3838 3886 3884 3898
rect 3838 3852 3844 3886
rect 3878 3852 3884 3886
rect 3838 3840 3884 3852
rect 3758 3258 3804 3270
rect 3758 3224 3764 3258
rect 3798 3224 3804 3258
rect 3758 3212 3804 3224
rect 3655 3014 3661 3066
rect 3713 3014 3719 3066
rect 672 3007 730 3013
rect 672 2973 684 3007
rect 718 2973 730 3007
rect 672 2967 730 2973
rect 592 2557 650 2563
rect 592 2523 604 2557
rect 638 2523 650 2557
rect 592 2517 650 2523
rect 3655 2464 3661 2516
rect 3713 2464 3719 2516
rect 3767 1690 3795 3212
rect 3847 2318 3875 3840
rect 3927 2480 3955 4002
rect 4007 3108 4035 4630
rect 3998 3096 4044 3108
rect 3998 3062 4004 3096
rect 4038 3062 4044 3096
rect 3998 3050 4044 3062
rect 3918 2468 3964 2480
rect 3918 2434 3924 2468
rect 3958 2434 3964 2468
rect 3918 2422 3964 2434
rect 3838 2306 3884 2318
rect 3838 2272 3844 2306
rect 3878 2272 3884 2306
rect 3838 2260 3884 2272
rect 3758 1678 3804 1690
rect 3758 1644 3764 1678
rect 3798 1644 3804 1678
rect 3758 1632 3804 1644
rect 3655 1434 3661 1486
rect 3713 1434 3719 1486
rect 3655 884 3661 936
rect 3713 884 3719 936
rect 3655 644 3661 696
rect 3713 644 3719 696
rect 672 637 730 643
rect 672 603 684 637
rect 718 603 730 637
rect 672 597 730 603
rect 3767 241 3795 1632
rect 3847 738 3875 2260
rect 3927 1031 3955 2422
rect 4007 1528 4035 3050
rect 4087 2402 4115 6484
rect 4167 2996 4195 8064
rect 4247 4576 4275 9644
rect 4327 6156 4355 11224
rect 4318 6144 4364 6156
rect 4318 6110 4324 6144
rect 4358 6110 4364 6144
rect 4318 6098 4364 6110
rect 4327 5752 4355 6098
rect 4407 6066 4435 25308
rect 4487 12386 4515 25308
rect 4567 18706 4595 25308
rect 4647 25026 4675 25308
rect 5023 25045 5029 25097
rect 5081 25045 5087 25097
rect 5495 25045 5501 25097
rect 5553 25045 5559 25097
rect 5927 25045 5933 25097
rect 5985 25045 5991 25097
rect 6271 25056 6277 25108
rect 6329 25056 6335 25108
rect 6695 25056 6701 25108
rect 6753 25056 6759 25108
rect 4638 25014 4684 25026
rect 4638 24980 4644 25014
rect 4678 24980 4684 25014
rect 4638 24968 4684 24980
rect 4647 24802 4675 24968
rect 4638 24790 4684 24802
rect 4638 24756 4644 24790
rect 4678 24756 4684 24790
rect 4638 24744 4684 24756
rect 4647 24236 4675 24744
rect 5023 24673 5029 24725
rect 5081 24673 5087 24725
rect 5495 24673 5501 24725
rect 5553 24673 5559 24725
rect 5927 24673 5933 24725
rect 5985 24673 5991 24725
rect 6271 24662 6277 24714
rect 6329 24662 6335 24714
rect 6695 24662 6701 24714
rect 6753 24662 6759 24714
rect 5023 24255 5029 24307
rect 5081 24255 5087 24307
rect 5495 24255 5501 24307
rect 5553 24255 5559 24307
rect 5927 24255 5933 24307
rect 5985 24255 5991 24307
rect 6271 24266 6277 24318
rect 6329 24266 6335 24318
rect 6695 24266 6701 24318
rect 6753 24266 6759 24318
rect 4638 24224 4684 24236
rect 4638 24190 4644 24224
rect 4678 24190 4684 24224
rect 4638 24178 4684 24190
rect 4647 24012 4675 24178
rect 4638 24000 4684 24012
rect 4638 23966 4644 24000
rect 4678 23966 4684 24000
rect 4638 23954 4684 23966
rect 4647 23446 4675 23954
rect 5023 23883 5029 23935
rect 5081 23883 5087 23935
rect 5495 23883 5501 23935
rect 5553 23883 5559 23935
rect 5927 23883 5933 23935
rect 5985 23883 5991 23935
rect 6271 23872 6277 23924
rect 6329 23872 6335 23924
rect 6695 23872 6701 23924
rect 6753 23872 6759 23924
rect 5023 23465 5029 23517
rect 5081 23465 5087 23517
rect 5495 23465 5501 23517
rect 5553 23465 5559 23517
rect 5927 23465 5933 23517
rect 5985 23465 5991 23517
rect 6271 23476 6277 23528
rect 6329 23476 6335 23528
rect 6695 23476 6701 23528
rect 6753 23476 6759 23528
rect 4638 23434 4684 23446
rect 4638 23400 4644 23434
rect 4678 23400 4684 23434
rect 4638 23388 4684 23400
rect 4647 23222 4675 23388
rect 4638 23210 4684 23222
rect 4638 23176 4644 23210
rect 4678 23176 4684 23210
rect 4638 23164 4684 23176
rect 4647 22656 4675 23164
rect 5023 23093 5029 23145
rect 5081 23093 5087 23145
rect 5495 23093 5501 23145
rect 5553 23093 5559 23145
rect 5927 23093 5933 23145
rect 5985 23093 5991 23145
rect 6271 23082 6277 23134
rect 6329 23082 6335 23134
rect 6695 23082 6701 23134
rect 6753 23082 6759 23134
rect 5023 22675 5029 22727
rect 5081 22675 5087 22727
rect 5495 22675 5501 22727
rect 5553 22675 5559 22727
rect 5927 22675 5933 22727
rect 5985 22675 5991 22727
rect 6271 22686 6277 22738
rect 6329 22686 6335 22738
rect 6695 22686 6701 22738
rect 6753 22686 6759 22738
rect 4638 22644 4684 22656
rect 4638 22610 4644 22644
rect 4678 22610 4684 22644
rect 4638 22598 4684 22610
rect 4647 22432 4675 22598
rect 4638 22420 4684 22432
rect 4638 22386 4644 22420
rect 4678 22386 4684 22420
rect 4638 22374 4684 22386
rect 4647 21866 4675 22374
rect 5023 22303 5029 22355
rect 5081 22303 5087 22355
rect 5495 22303 5501 22355
rect 5553 22303 5559 22355
rect 5927 22303 5933 22355
rect 5985 22303 5991 22355
rect 6271 22292 6277 22344
rect 6329 22292 6335 22344
rect 6695 22292 6701 22344
rect 6753 22292 6759 22344
rect 5023 21885 5029 21937
rect 5081 21885 5087 21937
rect 5495 21885 5501 21937
rect 5553 21885 5559 21937
rect 5927 21885 5933 21937
rect 5985 21885 5991 21937
rect 6271 21896 6277 21948
rect 6329 21896 6335 21948
rect 6695 21896 6701 21948
rect 6753 21896 6759 21948
rect 4638 21854 4684 21866
rect 4638 21820 4644 21854
rect 4678 21820 4684 21854
rect 4638 21808 4684 21820
rect 4647 21642 4675 21808
rect 4638 21630 4684 21642
rect 4638 21596 4644 21630
rect 4678 21596 4684 21630
rect 4638 21584 4684 21596
rect 4647 21076 4675 21584
rect 5023 21513 5029 21565
rect 5081 21513 5087 21565
rect 5495 21513 5501 21565
rect 5553 21513 5559 21565
rect 5927 21513 5933 21565
rect 5985 21513 5991 21565
rect 6271 21502 6277 21554
rect 6329 21502 6335 21554
rect 6695 21502 6701 21554
rect 6753 21502 6759 21554
rect 5023 21095 5029 21147
rect 5081 21095 5087 21147
rect 5495 21095 5501 21147
rect 5553 21095 5559 21147
rect 5927 21095 5933 21147
rect 5985 21095 5991 21147
rect 6271 21106 6277 21158
rect 6329 21106 6335 21158
rect 6695 21106 6701 21158
rect 6753 21106 6759 21158
rect 4638 21064 4684 21076
rect 4638 21030 4644 21064
rect 4678 21030 4684 21064
rect 4638 21018 4684 21030
rect 4647 20852 4675 21018
rect 4638 20840 4684 20852
rect 4638 20806 4644 20840
rect 4678 20806 4684 20840
rect 4638 20794 4684 20806
rect 4647 20286 4675 20794
rect 5023 20723 5029 20775
rect 5081 20723 5087 20775
rect 5495 20723 5501 20775
rect 5553 20723 5559 20775
rect 5927 20723 5933 20775
rect 5985 20723 5991 20775
rect 6271 20712 6277 20764
rect 6329 20712 6335 20764
rect 6695 20712 6701 20764
rect 6753 20712 6759 20764
rect 5023 20305 5029 20357
rect 5081 20305 5087 20357
rect 5495 20305 5501 20357
rect 5553 20305 5559 20357
rect 5927 20305 5933 20357
rect 5985 20305 5991 20357
rect 6271 20316 6277 20368
rect 6329 20316 6335 20368
rect 6695 20316 6701 20368
rect 6753 20316 6759 20368
rect 4638 20274 4684 20286
rect 4638 20240 4644 20274
rect 4678 20240 4684 20274
rect 4638 20228 4684 20240
rect 4647 20062 4675 20228
rect 4638 20050 4684 20062
rect 4638 20016 4644 20050
rect 4678 20016 4684 20050
rect 4638 20004 4684 20016
rect 4647 19496 4675 20004
rect 5023 19933 5029 19985
rect 5081 19933 5087 19985
rect 5495 19933 5501 19985
rect 5553 19933 5559 19985
rect 5927 19933 5933 19985
rect 5985 19933 5991 19985
rect 6271 19922 6277 19974
rect 6329 19922 6335 19974
rect 6695 19922 6701 19974
rect 6753 19922 6759 19974
rect 5023 19515 5029 19567
rect 5081 19515 5087 19567
rect 5495 19515 5501 19567
rect 5553 19515 5559 19567
rect 5927 19515 5933 19567
rect 5985 19515 5991 19567
rect 6271 19526 6277 19578
rect 6329 19526 6335 19578
rect 6695 19526 6701 19578
rect 6753 19526 6759 19578
rect 4638 19484 4684 19496
rect 4638 19450 4644 19484
rect 4678 19450 4684 19484
rect 4638 19438 4684 19450
rect 4647 19272 4675 19438
rect 4638 19260 4684 19272
rect 4638 19226 4644 19260
rect 4678 19226 4684 19260
rect 4638 19214 4684 19226
rect 4558 18694 4604 18706
rect 4558 18660 4564 18694
rect 4598 18660 4604 18694
rect 4558 18648 4604 18660
rect 4567 18482 4595 18648
rect 4558 18470 4604 18482
rect 4558 18436 4564 18470
rect 4598 18436 4604 18470
rect 4558 18424 4604 18436
rect 4567 17916 4595 18424
rect 4558 17904 4604 17916
rect 4558 17870 4564 17904
rect 4598 17870 4604 17904
rect 4558 17858 4604 17870
rect 4567 17692 4595 17858
rect 4558 17680 4604 17692
rect 4558 17646 4564 17680
rect 4598 17646 4604 17680
rect 4558 17634 4604 17646
rect 4567 17126 4595 17634
rect 4558 17114 4604 17126
rect 4558 17080 4564 17114
rect 4598 17080 4604 17114
rect 4558 17068 4604 17080
rect 4567 16902 4595 17068
rect 4558 16890 4604 16902
rect 4558 16856 4564 16890
rect 4598 16856 4604 16890
rect 4558 16844 4604 16856
rect 4567 16336 4595 16844
rect 4558 16324 4604 16336
rect 4558 16290 4564 16324
rect 4598 16290 4604 16324
rect 4558 16278 4604 16290
rect 4567 16112 4595 16278
rect 4558 16100 4604 16112
rect 4558 16066 4564 16100
rect 4598 16066 4604 16100
rect 4558 16054 4604 16066
rect 4567 15546 4595 16054
rect 4558 15534 4604 15546
rect 4558 15500 4564 15534
rect 4598 15500 4604 15534
rect 4558 15488 4604 15500
rect 4567 15322 4595 15488
rect 4558 15310 4604 15322
rect 4558 15276 4564 15310
rect 4598 15276 4604 15310
rect 4558 15264 4604 15276
rect 4567 14756 4595 15264
rect 4558 14744 4604 14756
rect 4558 14710 4564 14744
rect 4598 14710 4604 14744
rect 4558 14698 4604 14710
rect 4567 14532 4595 14698
rect 4558 14520 4604 14532
rect 4558 14486 4564 14520
rect 4598 14486 4604 14520
rect 4558 14474 4604 14486
rect 4567 13966 4595 14474
rect 4558 13954 4604 13966
rect 4558 13920 4564 13954
rect 4598 13920 4604 13954
rect 4558 13908 4604 13920
rect 4567 13742 4595 13908
rect 4558 13730 4604 13742
rect 4558 13696 4564 13730
rect 4598 13696 4604 13730
rect 4558 13684 4604 13696
rect 4567 13176 4595 13684
rect 4558 13164 4604 13176
rect 4558 13130 4564 13164
rect 4598 13130 4604 13164
rect 4558 13118 4604 13130
rect 4567 12952 4595 13118
rect 4558 12940 4604 12952
rect 4558 12906 4564 12940
rect 4598 12906 4604 12940
rect 4558 12894 4604 12906
rect 4478 12374 4524 12386
rect 4478 12340 4484 12374
rect 4518 12340 4524 12374
rect 4478 12328 4524 12340
rect 4487 12162 4515 12328
rect 4478 12150 4524 12162
rect 4478 12116 4484 12150
rect 4518 12116 4524 12150
rect 4478 12104 4524 12116
rect 4487 11596 4515 12104
rect 4478 11584 4524 11596
rect 4478 11550 4484 11584
rect 4518 11550 4524 11584
rect 4478 11538 4524 11550
rect 4487 11372 4515 11538
rect 4478 11360 4524 11372
rect 4478 11326 4484 11360
rect 4518 11326 4524 11360
rect 4478 11314 4524 11326
rect 4487 10806 4515 11314
rect 4478 10794 4524 10806
rect 4478 10760 4484 10794
rect 4518 10760 4524 10794
rect 4478 10748 4524 10760
rect 4487 10582 4515 10748
rect 4478 10570 4524 10582
rect 4478 10536 4484 10570
rect 4518 10536 4524 10570
rect 4478 10524 4524 10536
rect 4487 10016 4515 10524
rect 4478 10004 4524 10016
rect 4478 9970 4484 10004
rect 4518 9970 4524 10004
rect 4478 9958 4524 9970
rect 4487 9792 4515 9958
rect 4478 9780 4524 9792
rect 4478 9746 4484 9780
rect 4518 9746 4524 9780
rect 4478 9734 4524 9746
rect 4487 9226 4515 9734
rect 4478 9214 4524 9226
rect 4478 9180 4484 9214
rect 4518 9180 4524 9214
rect 4478 9168 4524 9180
rect 4487 9002 4515 9168
rect 4478 8990 4524 9002
rect 4478 8956 4484 8990
rect 4518 8956 4524 8990
rect 4478 8944 4524 8956
rect 4487 8436 4515 8944
rect 4478 8424 4524 8436
rect 4478 8390 4484 8424
rect 4518 8390 4524 8424
rect 4478 8378 4524 8390
rect 4487 8212 4515 8378
rect 4478 8200 4524 8212
rect 4478 8166 4484 8200
rect 4518 8166 4524 8200
rect 4478 8154 4524 8166
rect 4487 7646 4515 8154
rect 4478 7634 4524 7646
rect 4478 7600 4484 7634
rect 4518 7600 4524 7634
rect 4478 7588 4524 7600
rect 4487 7422 4515 7588
rect 4478 7410 4524 7422
rect 4478 7376 4484 7410
rect 4518 7376 4524 7410
rect 4478 7364 4524 7376
rect 4487 6856 4515 7364
rect 4478 6844 4524 6856
rect 4478 6810 4484 6844
rect 4518 6810 4524 6844
rect 4478 6798 4524 6810
rect 4487 6632 4515 6798
rect 4478 6620 4524 6632
rect 4478 6586 4484 6620
rect 4518 6586 4524 6620
rect 4478 6574 4524 6586
rect 4398 6054 4444 6066
rect 4398 6020 4404 6054
rect 4438 6020 4444 6054
rect 4398 6008 4444 6020
rect 4407 5842 4435 6008
rect 4398 5830 4444 5842
rect 4398 5796 4404 5830
rect 4438 5796 4444 5830
rect 4398 5784 4444 5796
rect 4318 5740 4364 5752
rect 4318 5706 4324 5740
rect 4358 5706 4364 5740
rect 4318 5694 4364 5706
rect 4327 5366 4355 5694
rect 4318 5354 4364 5366
rect 4318 5320 4324 5354
rect 4358 5320 4364 5354
rect 4318 5308 4364 5320
rect 4327 4962 4355 5308
rect 4407 5276 4435 5784
rect 4398 5264 4444 5276
rect 4398 5230 4404 5264
rect 4438 5230 4444 5264
rect 4398 5218 4444 5230
rect 4407 5052 4435 5218
rect 4487 5167 4515 6574
rect 4567 5562 4595 12894
rect 4647 5957 4675 19214
rect 5023 19143 5029 19195
rect 5081 19143 5087 19195
rect 5495 19143 5501 19195
rect 5553 19143 5559 19195
rect 5927 19143 5933 19195
rect 5985 19143 5991 19195
rect 6271 19132 6277 19184
rect 6329 19132 6335 19184
rect 6695 19132 6701 19184
rect 6753 19132 6759 19184
rect 5023 18725 5029 18777
rect 5081 18725 5087 18777
rect 5495 18725 5501 18777
rect 5553 18725 5559 18777
rect 5927 18725 5933 18777
rect 5985 18725 5991 18777
rect 6271 18736 6277 18788
rect 6329 18736 6335 18788
rect 6695 18736 6701 18788
rect 6753 18736 6759 18788
rect 5023 18353 5029 18405
rect 5081 18353 5087 18405
rect 5495 18353 5501 18405
rect 5553 18353 5559 18405
rect 5927 18353 5933 18405
rect 5985 18353 5991 18405
rect 6271 18342 6277 18394
rect 6329 18342 6335 18394
rect 6695 18342 6701 18394
rect 6753 18342 6759 18394
rect 5023 17935 5029 17987
rect 5081 17935 5087 17987
rect 5495 17935 5501 17987
rect 5553 17935 5559 17987
rect 5927 17935 5933 17987
rect 5985 17935 5991 17987
rect 6271 17946 6277 17998
rect 6329 17946 6335 17998
rect 6695 17946 6701 17998
rect 6753 17946 6759 17998
rect 5023 17563 5029 17615
rect 5081 17563 5087 17615
rect 5495 17563 5501 17615
rect 5553 17563 5559 17615
rect 5927 17563 5933 17615
rect 5985 17563 5991 17615
rect 6271 17552 6277 17604
rect 6329 17552 6335 17604
rect 6695 17552 6701 17604
rect 6753 17552 6759 17604
rect 5023 17145 5029 17197
rect 5081 17145 5087 17197
rect 5495 17145 5501 17197
rect 5553 17145 5559 17197
rect 5927 17145 5933 17197
rect 5985 17145 5991 17197
rect 6271 17156 6277 17208
rect 6329 17156 6335 17208
rect 6695 17156 6701 17208
rect 6753 17156 6759 17208
rect 5023 16773 5029 16825
rect 5081 16773 5087 16825
rect 5495 16773 5501 16825
rect 5553 16773 5559 16825
rect 5927 16773 5933 16825
rect 5985 16773 5991 16825
rect 6271 16762 6277 16814
rect 6329 16762 6335 16814
rect 6695 16762 6701 16814
rect 6753 16762 6759 16814
rect 5023 16355 5029 16407
rect 5081 16355 5087 16407
rect 5495 16355 5501 16407
rect 5553 16355 5559 16407
rect 5927 16355 5933 16407
rect 5985 16355 5991 16407
rect 6271 16366 6277 16418
rect 6329 16366 6335 16418
rect 6695 16366 6701 16418
rect 6753 16366 6759 16418
rect 5023 15983 5029 16035
rect 5081 15983 5087 16035
rect 5495 15983 5501 16035
rect 5553 15983 5559 16035
rect 5927 15983 5933 16035
rect 5985 15983 5991 16035
rect 6271 15972 6277 16024
rect 6329 15972 6335 16024
rect 6695 15972 6701 16024
rect 6753 15972 6759 16024
rect 5023 15565 5029 15617
rect 5081 15565 5087 15617
rect 5495 15565 5501 15617
rect 5553 15565 5559 15617
rect 5927 15565 5933 15617
rect 5985 15565 5991 15617
rect 6271 15576 6277 15628
rect 6329 15576 6335 15628
rect 6695 15576 6701 15628
rect 6753 15576 6759 15628
rect 5023 15193 5029 15245
rect 5081 15193 5087 15245
rect 5495 15193 5501 15245
rect 5553 15193 5559 15245
rect 5927 15193 5933 15245
rect 5985 15193 5991 15245
rect 6271 15182 6277 15234
rect 6329 15182 6335 15234
rect 6695 15182 6701 15234
rect 6753 15182 6759 15234
rect 5023 14775 5029 14827
rect 5081 14775 5087 14827
rect 5495 14775 5501 14827
rect 5553 14775 5559 14827
rect 5927 14775 5933 14827
rect 5985 14775 5991 14827
rect 6271 14786 6277 14838
rect 6329 14786 6335 14838
rect 6695 14786 6701 14838
rect 6753 14786 6759 14838
rect 5023 14403 5029 14455
rect 5081 14403 5087 14455
rect 5495 14403 5501 14455
rect 5553 14403 5559 14455
rect 5927 14403 5933 14455
rect 5985 14403 5991 14455
rect 6271 14392 6277 14444
rect 6329 14392 6335 14444
rect 6695 14392 6701 14444
rect 6753 14392 6759 14444
rect 5023 13985 5029 14037
rect 5081 13985 5087 14037
rect 5495 13985 5501 14037
rect 5553 13985 5559 14037
rect 5927 13985 5933 14037
rect 5985 13985 5991 14037
rect 6271 13996 6277 14048
rect 6329 13996 6335 14048
rect 6695 13996 6701 14048
rect 6753 13996 6759 14048
rect 5023 13613 5029 13665
rect 5081 13613 5087 13665
rect 5495 13613 5501 13665
rect 5553 13613 5559 13665
rect 5927 13613 5933 13665
rect 5985 13613 5991 13665
rect 6271 13602 6277 13654
rect 6329 13602 6335 13654
rect 6695 13602 6701 13654
rect 6753 13602 6759 13654
rect 5023 13195 5029 13247
rect 5081 13195 5087 13247
rect 5495 13195 5501 13247
rect 5553 13195 5559 13247
rect 5927 13195 5933 13247
rect 5985 13195 5991 13247
rect 6271 13206 6277 13258
rect 6329 13206 6335 13258
rect 6695 13206 6701 13258
rect 6753 13206 6759 13258
rect 5023 12823 5029 12875
rect 5081 12823 5087 12875
rect 5495 12823 5501 12875
rect 5553 12823 5559 12875
rect 5927 12823 5933 12875
rect 5985 12823 5991 12875
rect 6271 12812 6277 12864
rect 6329 12812 6335 12864
rect 6695 12812 6701 12864
rect 6753 12812 6759 12864
rect 5023 12405 5029 12457
rect 5081 12405 5087 12457
rect 5495 12405 5501 12457
rect 5553 12405 5559 12457
rect 5927 12405 5933 12457
rect 5985 12405 5991 12457
rect 6271 12416 6277 12468
rect 6329 12416 6335 12468
rect 6695 12416 6701 12468
rect 6753 12416 6759 12468
rect 5023 12033 5029 12085
rect 5081 12033 5087 12085
rect 5495 12033 5501 12085
rect 5553 12033 5559 12085
rect 5927 12033 5933 12085
rect 5985 12033 5991 12085
rect 6271 12022 6277 12074
rect 6329 12022 6335 12074
rect 6695 12022 6701 12074
rect 6753 12022 6759 12074
rect 5023 11615 5029 11667
rect 5081 11615 5087 11667
rect 5495 11615 5501 11667
rect 5553 11615 5559 11667
rect 5927 11615 5933 11667
rect 5985 11615 5991 11667
rect 6271 11626 6277 11678
rect 6329 11626 6335 11678
rect 6695 11626 6701 11678
rect 6753 11626 6759 11678
rect 5023 11243 5029 11295
rect 5081 11243 5087 11295
rect 5495 11243 5501 11295
rect 5553 11243 5559 11295
rect 5927 11243 5933 11295
rect 5985 11243 5991 11295
rect 6271 11232 6277 11284
rect 6329 11232 6335 11284
rect 6695 11232 6701 11284
rect 6753 11232 6759 11284
rect 5023 10825 5029 10877
rect 5081 10825 5087 10877
rect 5495 10825 5501 10877
rect 5553 10825 5559 10877
rect 5927 10825 5933 10877
rect 5985 10825 5991 10877
rect 6271 10836 6277 10888
rect 6329 10836 6335 10888
rect 6695 10836 6701 10888
rect 6753 10836 6759 10888
rect 5023 10453 5029 10505
rect 5081 10453 5087 10505
rect 5495 10453 5501 10505
rect 5553 10453 5559 10505
rect 5927 10453 5933 10505
rect 5985 10453 5991 10505
rect 6271 10442 6277 10494
rect 6329 10442 6335 10494
rect 6695 10442 6701 10494
rect 6753 10442 6759 10494
rect 5023 10035 5029 10087
rect 5081 10035 5087 10087
rect 5495 10035 5501 10087
rect 5553 10035 5559 10087
rect 5927 10035 5933 10087
rect 5985 10035 5991 10087
rect 6271 10046 6277 10098
rect 6329 10046 6335 10098
rect 6695 10046 6701 10098
rect 6753 10046 6759 10098
rect 5023 9663 5029 9715
rect 5081 9663 5087 9715
rect 5495 9663 5501 9715
rect 5553 9663 5559 9715
rect 5927 9663 5933 9715
rect 5985 9663 5991 9715
rect 6271 9652 6277 9704
rect 6329 9652 6335 9704
rect 6695 9652 6701 9704
rect 6753 9652 6759 9704
rect 5023 9245 5029 9297
rect 5081 9245 5087 9297
rect 5495 9245 5501 9297
rect 5553 9245 5559 9297
rect 5927 9245 5933 9297
rect 5985 9245 5991 9297
rect 6271 9256 6277 9308
rect 6329 9256 6335 9308
rect 6695 9256 6701 9308
rect 6753 9256 6759 9308
rect 5023 8873 5029 8925
rect 5081 8873 5087 8925
rect 5495 8873 5501 8925
rect 5553 8873 5559 8925
rect 5927 8873 5933 8925
rect 5985 8873 5991 8925
rect 6271 8862 6277 8914
rect 6329 8862 6335 8914
rect 6695 8862 6701 8914
rect 6753 8862 6759 8914
rect 5023 8455 5029 8507
rect 5081 8455 5087 8507
rect 5495 8455 5501 8507
rect 5553 8455 5559 8507
rect 5927 8455 5933 8507
rect 5985 8455 5991 8507
rect 6271 8466 6277 8518
rect 6329 8466 6335 8518
rect 6695 8466 6701 8518
rect 6753 8466 6759 8518
rect 5023 8083 5029 8135
rect 5081 8083 5087 8135
rect 5495 8083 5501 8135
rect 5553 8083 5559 8135
rect 5927 8083 5933 8135
rect 5985 8083 5991 8135
rect 6271 8072 6277 8124
rect 6329 8072 6335 8124
rect 6695 8072 6701 8124
rect 6753 8072 6759 8124
rect 5023 7665 5029 7717
rect 5081 7665 5087 7717
rect 5495 7665 5501 7717
rect 5553 7665 5559 7717
rect 5927 7665 5933 7717
rect 5985 7665 5991 7717
rect 6271 7676 6277 7728
rect 6329 7676 6335 7728
rect 6695 7676 6701 7728
rect 6753 7676 6759 7728
rect 5023 7293 5029 7345
rect 5081 7293 5087 7345
rect 5495 7293 5501 7345
rect 5553 7293 5559 7345
rect 5927 7293 5933 7345
rect 5985 7293 5991 7345
rect 6271 7282 6277 7334
rect 6329 7282 6335 7334
rect 6695 7282 6701 7334
rect 6753 7282 6759 7334
rect 5023 6875 5029 6927
rect 5081 6875 5087 6927
rect 5495 6875 5501 6927
rect 5553 6875 5559 6927
rect 5927 6875 5933 6927
rect 5985 6875 5991 6927
rect 6271 6886 6277 6938
rect 6329 6886 6335 6938
rect 6695 6886 6701 6938
rect 6753 6886 6759 6938
rect 5023 6503 5029 6555
rect 5081 6503 5087 6555
rect 5495 6503 5501 6555
rect 5553 6503 5559 6555
rect 5927 6503 5933 6555
rect 5985 6503 5991 6555
rect 6271 6492 6277 6544
rect 6329 6492 6335 6544
rect 6695 6492 6701 6544
rect 6753 6492 6759 6544
rect 5023 6085 5029 6137
rect 5081 6085 5087 6137
rect 5495 6085 5501 6137
rect 5553 6085 5559 6137
rect 5927 6085 5933 6137
rect 5985 6085 5991 6137
rect 6271 6096 6277 6148
rect 6329 6096 6335 6148
rect 6695 6096 6701 6148
rect 6753 6096 6759 6148
rect 4635 5951 4687 5957
rect 4635 5893 4687 5899
rect 4555 5556 4607 5562
rect 4555 5498 4607 5504
rect 4475 5161 4527 5167
rect 4475 5103 4527 5109
rect 4398 5040 4444 5052
rect 4398 5006 4404 5040
rect 4438 5006 4444 5040
rect 4398 4994 4444 5006
rect 4318 4950 4364 4962
rect 4318 4916 4324 4950
rect 4358 4916 4364 4950
rect 4318 4904 4364 4916
rect 4238 4564 4284 4576
rect 4238 4530 4244 4564
rect 4278 4530 4284 4564
rect 4238 4518 4284 4530
rect 4247 4172 4275 4518
rect 4238 4160 4284 4172
rect 4238 4126 4244 4160
rect 4278 4126 4284 4160
rect 4238 4114 4284 4126
rect 4247 3786 4275 4114
rect 4238 3774 4284 3786
rect 4238 3740 4244 3774
rect 4278 3740 4284 3774
rect 4238 3728 4284 3740
rect 4247 3382 4275 3728
rect 4327 3587 4355 4904
rect 4407 4772 4435 4994
rect 4395 4766 4447 4772
rect 4395 4708 4447 4714
rect 4407 4486 4435 4708
rect 4398 4474 4444 4486
rect 4398 4440 4404 4474
rect 4438 4440 4444 4474
rect 4398 4428 4444 4440
rect 4407 4262 4435 4428
rect 4398 4250 4444 4262
rect 4398 4216 4404 4250
rect 4438 4216 4444 4250
rect 4398 4204 4444 4216
rect 4407 3696 4435 4204
rect 4398 3684 4444 3696
rect 4398 3650 4404 3684
rect 4438 3650 4444 3684
rect 4398 3638 4444 3650
rect 4315 3581 4367 3587
rect 4315 3523 4367 3529
rect 4238 3370 4284 3382
rect 4238 3336 4244 3370
rect 4278 3336 4284 3370
rect 4238 3324 4284 3336
rect 4247 3192 4275 3324
rect 4235 3186 4287 3192
rect 4235 3128 4287 3134
rect 4158 2984 4204 2996
rect 4158 2950 4164 2984
rect 4198 2950 4204 2984
rect 4158 2938 4204 2950
rect 4167 2797 4195 2938
rect 4155 2791 4207 2797
rect 4155 2733 4207 2739
rect 4167 2592 4195 2733
rect 4158 2580 4204 2592
rect 4158 2546 4164 2580
rect 4198 2546 4204 2580
rect 4158 2534 4204 2546
rect 4075 2396 4127 2402
rect 4075 2338 4127 2344
rect 3998 1516 4044 1528
rect 3998 1482 4004 1516
rect 4038 1482 4044 1516
rect 3998 1470 4044 1482
rect 4007 1217 4035 1470
rect 4087 1416 4115 2338
rect 4167 2206 4195 2534
rect 4158 2194 4204 2206
rect 4158 2160 4164 2194
rect 4198 2160 4204 2194
rect 4158 2148 4204 2160
rect 4167 1802 4195 2148
rect 4158 1790 4204 1802
rect 4158 1756 4164 1790
rect 4198 1756 4204 1790
rect 4158 1744 4204 1756
rect 4078 1404 4124 1416
rect 4078 1370 4084 1404
rect 4118 1370 4124 1404
rect 4078 1358 4124 1370
rect 3995 1211 4047 1217
rect 3995 1153 4047 1159
rect 3915 1025 3967 1031
rect 3915 967 3967 973
rect 3927 900 3955 967
rect 3918 888 3964 900
rect 3918 854 3924 888
rect 3958 854 3964 888
rect 3918 842 3964 854
rect 3838 726 3884 738
rect 3838 692 3844 726
rect 3878 692 3884 726
rect 3838 680 3884 692
rect 3847 427 3875 680
rect 3835 421 3887 427
rect 3835 363 3887 369
rect 3755 235 3807 241
rect 592 187 650 193
rect 592 153 604 187
rect 638 153 650 187
rect 3755 177 3807 183
rect 592 147 650 153
rect 3655 94 3661 146
rect 3713 94 3719 146
rect 3767 110 3795 177
rect 3758 98 3804 110
rect 3758 64 3764 98
rect 3798 64 3804 98
rect 3758 52 3804 64
rect 3767 0 3795 52
rect 3847 0 3875 363
rect 3927 0 3955 842
rect 4007 0 4035 1153
rect 4087 1012 4115 1358
rect 4078 1000 4124 1012
rect 4078 966 4084 1000
rect 4118 966 4124 1000
rect 4078 954 4124 966
rect 4087 626 4115 954
rect 4078 614 4124 626
rect 4078 580 4084 614
rect 4118 580 4124 614
rect 4078 568 4124 580
rect 4087 222 4115 568
rect 4078 210 4124 222
rect 4078 176 4084 210
rect 4118 176 4124 210
rect 4078 164 4124 176
rect 4087 0 4115 164
rect 4167 0 4195 1744
rect 4247 0 4275 3128
rect 4327 0 4355 3523
rect 4407 3472 4435 3638
rect 4398 3460 4444 3472
rect 4398 3426 4404 3460
rect 4438 3426 4444 3460
rect 4398 3414 4444 3426
rect 4407 2906 4435 3414
rect 4398 2894 4444 2906
rect 4398 2860 4404 2894
rect 4438 2860 4444 2894
rect 4398 2848 4444 2860
rect 4407 2682 4435 2848
rect 4398 2670 4444 2682
rect 4398 2636 4404 2670
rect 4438 2636 4444 2670
rect 4398 2624 4444 2636
rect 4407 2116 4435 2624
rect 4398 2104 4444 2116
rect 4398 2070 4404 2104
rect 4438 2070 4444 2104
rect 4398 2058 4444 2070
rect 4407 1892 4435 2058
rect 4398 1880 4444 1892
rect 4398 1846 4404 1880
rect 4438 1846 4444 1880
rect 4398 1834 4444 1846
rect 4407 1326 4435 1834
rect 4398 1314 4444 1326
rect 4398 1280 4404 1314
rect 4438 1280 4444 1314
rect 4398 1268 4444 1280
rect 4407 1102 4435 1268
rect 4398 1090 4444 1102
rect 4398 1056 4404 1090
rect 4438 1056 4444 1090
rect 4398 1044 4444 1056
rect 4407 536 4435 1044
rect 4398 524 4444 536
rect 4398 490 4404 524
rect 4438 490 4444 524
rect 4398 478 4444 490
rect 4407 312 4435 478
rect 4398 300 4444 312
rect 4398 266 4404 300
rect 4438 266 4444 300
rect 4398 254 4444 266
rect 4407 0 4435 254
rect 4487 0 4515 5103
rect 4567 0 4595 5498
rect 4647 0 4675 5893
rect 5023 5713 5029 5765
rect 5081 5713 5087 5765
rect 5495 5713 5501 5765
rect 5553 5713 5559 5765
rect 5927 5713 5933 5765
rect 5985 5713 5991 5765
rect 6271 5702 6277 5754
rect 6329 5702 6335 5754
rect 6695 5702 6701 5754
rect 6753 5702 6759 5754
rect 5023 5295 5029 5347
rect 5081 5295 5087 5347
rect 5495 5295 5501 5347
rect 5553 5295 5559 5347
rect 5927 5295 5933 5347
rect 5985 5295 5991 5347
rect 6271 5306 6277 5358
rect 6329 5306 6335 5358
rect 6695 5306 6701 5358
rect 6753 5306 6759 5358
rect 5023 4923 5029 4975
rect 5081 4923 5087 4975
rect 5495 4923 5501 4975
rect 5553 4923 5559 4975
rect 5927 4923 5933 4975
rect 5985 4923 5991 4975
rect 6271 4912 6277 4964
rect 6329 4912 6335 4964
rect 6695 4912 6701 4964
rect 6753 4912 6759 4964
rect 5023 4505 5029 4557
rect 5081 4505 5087 4557
rect 5495 4505 5501 4557
rect 5553 4505 5559 4557
rect 5927 4505 5933 4557
rect 5985 4505 5991 4557
rect 6271 4516 6277 4568
rect 6329 4516 6335 4568
rect 6695 4516 6701 4568
rect 6753 4516 6759 4568
rect 5023 4133 5029 4185
rect 5081 4133 5087 4185
rect 5495 4133 5501 4185
rect 5553 4133 5559 4185
rect 5927 4133 5933 4185
rect 5985 4133 5991 4185
rect 6271 4122 6277 4174
rect 6329 4122 6335 4174
rect 6695 4122 6701 4174
rect 6753 4122 6759 4174
rect 5023 3715 5029 3767
rect 5081 3715 5087 3767
rect 5495 3715 5501 3767
rect 5553 3715 5559 3767
rect 5927 3715 5933 3767
rect 5985 3715 5991 3767
rect 6271 3726 6277 3778
rect 6329 3726 6335 3778
rect 6695 3726 6701 3778
rect 6753 3726 6759 3778
rect 5023 3343 5029 3395
rect 5081 3343 5087 3395
rect 5495 3343 5501 3395
rect 5553 3343 5559 3395
rect 5927 3343 5933 3395
rect 5985 3343 5991 3395
rect 6271 3332 6277 3384
rect 6329 3332 6335 3384
rect 6695 3332 6701 3384
rect 6753 3332 6759 3384
rect 5023 2925 5029 2977
rect 5081 2925 5087 2977
rect 5495 2925 5501 2977
rect 5553 2925 5559 2977
rect 5927 2925 5933 2977
rect 5985 2925 5991 2977
rect 6271 2936 6277 2988
rect 6329 2936 6335 2988
rect 6695 2936 6701 2988
rect 6753 2936 6759 2988
rect 5023 2553 5029 2605
rect 5081 2553 5087 2605
rect 5495 2553 5501 2605
rect 5553 2553 5559 2605
rect 5927 2553 5933 2605
rect 5985 2553 5991 2605
rect 6271 2542 6277 2594
rect 6329 2542 6335 2594
rect 6695 2542 6701 2594
rect 6753 2542 6759 2594
rect 5023 2135 5029 2187
rect 5081 2135 5087 2187
rect 5495 2135 5501 2187
rect 5553 2135 5559 2187
rect 5927 2135 5933 2187
rect 5985 2135 5991 2187
rect 6271 2146 6277 2198
rect 6329 2146 6335 2198
rect 6695 2146 6701 2198
rect 6753 2146 6759 2198
rect 5023 1763 5029 1815
rect 5081 1763 5087 1815
rect 5495 1763 5501 1815
rect 5553 1763 5559 1815
rect 5927 1763 5933 1815
rect 5985 1763 5991 1815
rect 6271 1752 6277 1804
rect 6329 1752 6335 1804
rect 6695 1752 6701 1804
rect 6753 1752 6759 1804
rect 5023 1345 5029 1397
rect 5081 1345 5087 1397
rect 5495 1345 5501 1397
rect 5553 1345 5559 1397
rect 5927 1345 5933 1397
rect 5985 1345 5991 1397
rect 6271 1356 6277 1408
rect 6329 1356 6335 1408
rect 6695 1356 6701 1408
rect 6753 1356 6759 1408
rect 5023 973 5029 1025
rect 5081 973 5087 1025
rect 5495 973 5501 1025
rect 5553 973 5559 1025
rect 5927 973 5933 1025
rect 5985 973 5991 1025
rect 6271 962 6277 1014
rect 6329 962 6335 1014
rect 6695 962 6701 1014
rect 6753 962 6759 1014
rect 5023 555 5029 607
rect 5081 555 5087 607
rect 5495 555 5501 607
rect 5553 555 5559 607
rect 5927 555 5933 607
rect 5985 555 5991 607
rect 6271 566 6277 618
rect 6329 566 6335 618
rect 6695 566 6701 618
rect 6753 566 6759 618
rect 5023 183 5029 235
rect 5081 183 5087 235
rect 5495 183 5501 235
rect 5553 183 5559 235
rect 5927 183 5933 235
rect 5985 183 5991 235
rect 6271 172 6277 224
rect 6329 172 6335 224
rect 6695 172 6701 224
rect 6753 172 6759 224
<< via1 >>
rect 3661 6217 3713 6226
rect 3661 6183 3670 6217
rect 3670 6183 3704 6217
rect 3704 6183 3713 6217
rect 3661 6174 3713 6183
rect 3661 5667 3713 5676
rect 3661 5633 3670 5667
rect 3670 5633 3704 5667
rect 3704 5633 3713 5667
rect 3661 5624 3713 5633
rect 3661 5427 3713 5436
rect 3661 5393 3670 5427
rect 3670 5393 3704 5427
rect 3704 5393 3713 5427
rect 3661 5384 3713 5393
rect 3661 4877 3713 4886
rect 3661 4843 3670 4877
rect 3670 4843 3704 4877
rect 3704 4843 3713 4877
rect 3661 4834 3713 4843
rect 3661 3847 3713 3856
rect 3661 3813 3670 3847
rect 3670 3813 3704 3847
rect 3704 3813 3713 3847
rect 3661 3804 3713 3813
rect 3661 3297 3713 3306
rect 3661 3263 3670 3297
rect 3670 3263 3704 3297
rect 3704 3263 3713 3297
rect 3661 3254 3713 3263
rect 3661 3057 3713 3066
rect 3661 3023 3670 3057
rect 3670 3023 3704 3057
rect 3704 3023 3713 3057
rect 3661 3014 3713 3023
rect 3661 2507 3713 2516
rect 3661 2473 3670 2507
rect 3670 2473 3704 2507
rect 3704 2473 3713 2507
rect 3661 2464 3713 2473
rect 3661 1477 3713 1486
rect 3661 1443 3670 1477
rect 3670 1443 3704 1477
rect 3704 1443 3713 1477
rect 3661 1434 3713 1443
rect 3661 927 3713 936
rect 3661 893 3670 927
rect 3670 893 3704 927
rect 3704 893 3713 927
rect 3661 884 3713 893
rect 3661 687 3713 696
rect 3661 653 3670 687
rect 3670 653 3704 687
rect 3704 653 3713 687
rect 3661 644 3713 653
rect 5029 25045 5081 25097
rect 5501 25045 5553 25097
rect 5933 25045 5985 25097
rect 6277 25056 6329 25108
rect 6701 25056 6753 25108
rect 5029 24673 5081 24725
rect 5501 24673 5553 24725
rect 5933 24673 5985 24725
rect 6277 24662 6329 24714
rect 6701 24662 6753 24714
rect 5029 24255 5081 24307
rect 5501 24255 5553 24307
rect 5933 24255 5985 24307
rect 6277 24266 6329 24318
rect 6701 24266 6753 24318
rect 5029 23883 5081 23935
rect 5501 23883 5553 23935
rect 5933 23883 5985 23935
rect 6277 23872 6329 23924
rect 6701 23872 6753 23924
rect 5029 23465 5081 23517
rect 5501 23465 5553 23517
rect 5933 23465 5985 23517
rect 6277 23476 6329 23528
rect 6701 23476 6753 23528
rect 5029 23093 5081 23145
rect 5501 23093 5553 23145
rect 5933 23093 5985 23145
rect 6277 23082 6329 23134
rect 6701 23082 6753 23134
rect 5029 22675 5081 22727
rect 5501 22675 5553 22727
rect 5933 22675 5985 22727
rect 6277 22686 6329 22738
rect 6701 22686 6753 22738
rect 5029 22303 5081 22355
rect 5501 22303 5553 22355
rect 5933 22303 5985 22355
rect 6277 22292 6329 22344
rect 6701 22292 6753 22344
rect 5029 21885 5081 21937
rect 5501 21885 5553 21937
rect 5933 21885 5985 21937
rect 6277 21896 6329 21948
rect 6701 21896 6753 21948
rect 5029 21513 5081 21565
rect 5501 21513 5553 21565
rect 5933 21513 5985 21565
rect 6277 21502 6329 21554
rect 6701 21502 6753 21554
rect 5029 21095 5081 21147
rect 5501 21095 5553 21147
rect 5933 21095 5985 21147
rect 6277 21106 6329 21158
rect 6701 21106 6753 21158
rect 5029 20723 5081 20775
rect 5501 20723 5553 20775
rect 5933 20723 5985 20775
rect 6277 20712 6329 20764
rect 6701 20712 6753 20764
rect 5029 20305 5081 20357
rect 5501 20305 5553 20357
rect 5933 20305 5985 20357
rect 6277 20316 6329 20368
rect 6701 20316 6753 20368
rect 5029 19933 5081 19985
rect 5501 19933 5553 19985
rect 5933 19933 5985 19985
rect 6277 19922 6329 19974
rect 6701 19922 6753 19974
rect 5029 19515 5081 19567
rect 5501 19515 5553 19567
rect 5933 19515 5985 19567
rect 6277 19526 6329 19578
rect 6701 19526 6753 19578
rect 5029 19143 5081 19195
rect 5501 19143 5553 19195
rect 5933 19143 5985 19195
rect 6277 19132 6329 19184
rect 6701 19132 6753 19184
rect 5029 18725 5081 18777
rect 5501 18725 5553 18777
rect 5933 18725 5985 18777
rect 6277 18736 6329 18788
rect 6701 18736 6753 18788
rect 5029 18353 5081 18405
rect 5501 18353 5553 18405
rect 5933 18353 5985 18405
rect 6277 18342 6329 18394
rect 6701 18342 6753 18394
rect 5029 17935 5081 17987
rect 5501 17935 5553 17987
rect 5933 17935 5985 17987
rect 6277 17946 6329 17998
rect 6701 17946 6753 17998
rect 5029 17563 5081 17615
rect 5501 17563 5553 17615
rect 5933 17563 5985 17615
rect 6277 17552 6329 17604
rect 6701 17552 6753 17604
rect 5029 17145 5081 17197
rect 5501 17145 5553 17197
rect 5933 17145 5985 17197
rect 6277 17156 6329 17208
rect 6701 17156 6753 17208
rect 5029 16773 5081 16825
rect 5501 16773 5553 16825
rect 5933 16773 5985 16825
rect 6277 16762 6329 16814
rect 6701 16762 6753 16814
rect 5029 16355 5081 16407
rect 5501 16355 5553 16407
rect 5933 16355 5985 16407
rect 6277 16366 6329 16418
rect 6701 16366 6753 16418
rect 5029 15983 5081 16035
rect 5501 15983 5553 16035
rect 5933 15983 5985 16035
rect 6277 15972 6329 16024
rect 6701 15972 6753 16024
rect 5029 15565 5081 15617
rect 5501 15565 5553 15617
rect 5933 15565 5985 15617
rect 6277 15576 6329 15628
rect 6701 15576 6753 15628
rect 5029 15193 5081 15245
rect 5501 15193 5553 15245
rect 5933 15193 5985 15245
rect 6277 15182 6329 15234
rect 6701 15182 6753 15234
rect 5029 14775 5081 14827
rect 5501 14775 5553 14827
rect 5933 14775 5985 14827
rect 6277 14786 6329 14838
rect 6701 14786 6753 14838
rect 5029 14403 5081 14455
rect 5501 14403 5553 14455
rect 5933 14403 5985 14455
rect 6277 14392 6329 14444
rect 6701 14392 6753 14444
rect 5029 13985 5081 14037
rect 5501 13985 5553 14037
rect 5933 13985 5985 14037
rect 6277 13996 6329 14048
rect 6701 13996 6753 14048
rect 5029 13613 5081 13665
rect 5501 13613 5553 13665
rect 5933 13613 5985 13665
rect 6277 13602 6329 13654
rect 6701 13602 6753 13654
rect 5029 13195 5081 13247
rect 5501 13195 5553 13247
rect 5933 13195 5985 13247
rect 6277 13206 6329 13258
rect 6701 13206 6753 13258
rect 5029 12823 5081 12875
rect 5501 12823 5553 12875
rect 5933 12823 5985 12875
rect 6277 12812 6329 12864
rect 6701 12812 6753 12864
rect 5029 12405 5081 12457
rect 5501 12405 5553 12457
rect 5933 12405 5985 12457
rect 6277 12416 6329 12468
rect 6701 12416 6753 12468
rect 5029 12033 5081 12085
rect 5501 12033 5553 12085
rect 5933 12033 5985 12085
rect 6277 12022 6329 12074
rect 6701 12022 6753 12074
rect 5029 11615 5081 11667
rect 5501 11615 5553 11667
rect 5933 11615 5985 11667
rect 6277 11626 6329 11678
rect 6701 11626 6753 11678
rect 5029 11243 5081 11295
rect 5501 11243 5553 11295
rect 5933 11243 5985 11295
rect 6277 11232 6329 11284
rect 6701 11232 6753 11284
rect 5029 10825 5081 10877
rect 5501 10825 5553 10877
rect 5933 10825 5985 10877
rect 6277 10836 6329 10888
rect 6701 10836 6753 10888
rect 5029 10453 5081 10505
rect 5501 10453 5553 10505
rect 5933 10453 5985 10505
rect 6277 10442 6329 10494
rect 6701 10442 6753 10494
rect 5029 10035 5081 10087
rect 5501 10035 5553 10087
rect 5933 10035 5985 10087
rect 6277 10046 6329 10098
rect 6701 10046 6753 10098
rect 5029 9663 5081 9715
rect 5501 9663 5553 9715
rect 5933 9663 5985 9715
rect 6277 9652 6329 9704
rect 6701 9652 6753 9704
rect 5029 9245 5081 9297
rect 5501 9245 5553 9297
rect 5933 9245 5985 9297
rect 6277 9256 6329 9308
rect 6701 9256 6753 9308
rect 5029 8873 5081 8925
rect 5501 8873 5553 8925
rect 5933 8873 5985 8925
rect 6277 8862 6329 8914
rect 6701 8862 6753 8914
rect 5029 8455 5081 8507
rect 5501 8455 5553 8507
rect 5933 8455 5985 8507
rect 6277 8466 6329 8518
rect 6701 8466 6753 8518
rect 5029 8083 5081 8135
rect 5501 8083 5553 8135
rect 5933 8083 5985 8135
rect 6277 8072 6329 8124
rect 6701 8072 6753 8124
rect 5029 7665 5081 7717
rect 5501 7665 5553 7717
rect 5933 7665 5985 7717
rect 6277 7676 6329 7728
rect 6701 7676 6753 7728
rect 5029 7293 5081 7345
rect 5501 7293 5553 7345
rect 5933 7293 5985 7345
rect 6277 7282 6329 7334
rect 6701 7282 6753 7334
rect 5029 6875 5081 6927
rect 5501 6875 5553 6927
rect 5933 6875 5985 6927
rect 6277 6886 6329 6938
rect 6701 6886 6753 6938
rect 5029 6503 5081 6555
rect 5501 6503 5553 6555
rect 5933 6503 5985 6555
rect 6277 6492 6329 6544
rect 6701 6492 6753 6544
rect 5029 6085 5081 6137
rect 5501 6085 5553 6137
rect 5933 6085 5985 6137
rect 6277 6096 6329 6148
rect 6701 6096 6753 6148
rect 4635 5899 4687 5951
rect 4555 5504 4607 5556
rect 4475 5109 4527 5161
rect 4395 4714 4447 4766
rect 4315 3529 4367 3581
rect 4235 3134 4287 3186
rect 4155 2739 4207 2791
rect 4075 2344 4127 2396
rect 3995 1159 4047 1211
rect 3915 973 3967 1025
rect 3835 369 3887 421
rect 3755 183 3807 235
rect 3661 137 3713 146
rect 3661 103 3670 137
rect 3670 103 3704 137
rect 3704 103 3713 137
rect 3661 94 3713 103
rect 5029 5713 5081 5765
rect 5501 5713 5553 5765
rect 5933 5713 5985 5765
rect 6277 5702 6329 5754
rect 6701 5702 6753 5754
rect 5029 5295 5081 5347
rect 5501 5295 5553 5347
rect 5933 5295 5985 5347
rect 6277 5306 6329 5358
rect 6701 5306 6753 5358
rect 5029 4923 5081 4975
rect 5501 4923 5553 4975
rect 5933 4923 5985 4975
rect 6277 4912 6329 4964
rect 6701 4912 6753 4964
rect 5029 4505 5081 4557
rect 5501 4505 5553 4557
rect 5933 4505 5985 4557
rect 6277 4516 6329 4568
rect 6701 4516 6753 4568
rect 5029 4133 5081 4185
rect 5501 4133 5553 4185
rect 5933 4133 5985 4185
rect 6277 4122 6329 4174
rect 6701 4122 6753 4174
rect 5029 3715 5081 3767
rect 5501 3715 5553 3767
rect 5933 3715 5985 3767
rect 6277 3726 6329 3778
rect 6701 3726 6753 3778
rect 5029 3343 5081 3395
rect 5501 3343 5553 3395
rect 5933 3343 5985 3395
rect 6277 3332 6329 3384
rect 6701 3332 6753 3384
rect 5029 2925 5081 2977
rect 5501 2925 5553 2977
rect 5933 2925 5985 2977
rect 6277 2936 6329 2988
rect 6701 2936 6753 2988
rect 5029 2553 5081 2605
rect 5501 2553 5553 2605
rect 5933 2553 5985 2605
rect 6277 2542 6329 2594
rect 6701 2542 6753 2594
rect 5029 2135 5081 2187
rect 5501 2135 5553 2187
rect 5933 2135 5985 2187
rect 6277 2146 6329 2198
rect 6701 2146 6753 2198
rect 5029 1763 5081 1815
rect 5501 1763 5553 1815
rect 5933 1763 5985 1815
rect 6277 1752 6329 1804
rect 6701 1752 6753 1804
rect 5029 1345 5081 1397
rect 5501 1345 5553 1397
rect 5933 1345 5985 1397
rect 6277 1356 6329 1408
rect 6701 1356 6753 1408
rect 5029 973 5081 1025
rect 5501 973 5553 1025
rect 5933 973 5985 1025
rect 6277 962 6329 1014
rect 6701 962 6753 1014
rect 5029 555 5081 607
rect 5501 555 5553 607
rect 5933 555 5985 607
rect 6277 566 6329 618
rect 6701 566 6753 618
rect 5029 183 5081 235
rect 5501 183 5553 235
rect 5933 183 5985 235
rect 6277 172 6329 224
rect 6701 172 6753 224
<< metal2 >>
rect 6275 25111 6331 25120
rect 5027 25099 5083 25108
rect 5027 25034 5083 25043
rect 5499 25099 5555 25108
rect 5499 25034 5555 25043
rect 5931 25099 5987 25108
rect 6275 25046 6331 25055
rect 6699 25111 6755 25120
rect 6699 25046 6755 25055
rect 5931 25034 5987 25043
rect 5027 24727 5083 24736
rect 5027 24662 5083 24671
rect 5499 24727 5555 24736
rect 5499 24662 5555 24671
rect 5931 24727 5987 24736
rect 5931 24662 5987 24671
rect 6275 24715 6331 24724
rect 6275 24650 6331 24659
rect 6699 24715 6755 24724
rect 6699 24650 6755 24659
rect 6275 24321 6331 24330
rect 5027 24309 5083 24318
rect 5027 24244 5083 24253
rect 5499 24309 5555 24318
rect 5499 24244 5555 24253
rect 5931 24309 5987 24318
rect 6275 24256 6331 24265
rect 6699 24321 6755 24330
rect 6699 24256 6755 24265
rect 5931 24244 5987 24253
rect 5027 23937 5083 23946
rect 5027 23872 5083 23881
rect 5499 23937 5555 23946
rect 5499 23872 5555 23881
rect 5931 23937 5987 23946
rect 5931 23872 5987 23881
rect 6275 23925 6331 23934
rect 6275 23860 6331 23869
rect 6699 23925 6755 23934
rect 6699 23860 6755 23869
rect 6275 23531 6331 23540
rect 5027 23519 5083 23528
rect 5027 23454 5083 23463
rect 5499 23519 5555 23528
rect 5499 23454 5555 23463
rect 5931 23519 5987 23528
rect 6275 23466 6331 23475
rect 6699 23531 6755 23540
rect 6699 23466 6755 23475
rect 5931 23454 5987 23463
rect 5027 23147 5083 23156
rect 5027 23082 5083 23091
rect 5499 23147 5555 23156
rect 5499 23082 5555 23091
rect 5931 23147 5987 23156
rect 5931 23082 5987 23091
rect 6275 23135 6331 23144
rect 6275 23070 6331 23079
rect 6699 23135 6755 23144
rect 6699 23070 6755 23079
rect 6275 22741 6331 22750
rect 5027 22729 5083 22738
rect 5027 22664 5083 22673
rect 5499 22729 5555 22738
rect 5499 22664 5555 22673
rect 5931 22729 5987 22738
rect 6275 22676 6331 22685
rect 6699 22741 6755 22750
rect 6699 22676 6755 22685
rect 5931 22664 5987 22673
rect 5027 22357 5083 22366
rect 5027 22292 5083 22301
rect 5499 22357 5555 22366
rect 5499 22292 5555 22301
rect 5931 22357 5987 22366
rect 5931 22292 5987 22301
rect 6275 22345 6331 22354
rect 6275 22280 6331 22289
rect 6699 22345 6755 22354
rect 6699 22280 6755 22289
rect 6275 21951 6331 21960
rect 5027 21939 5083 21948
rect 5027 21874 5083 21883
rect 5499 21939 5555 21948
rect 5499 21874 5555 21883
rect 5931 21939 5987 21948
rect 6275 21886 6331 21895
rect 6699 21951 6755 21960
rect 6699 21886 6755 21895
rect 5931 21874 5987 21883
rect 5027 21567 5083 21576
rect 5027 21502 5083 21511
rect 5499 21567 5555 21576
rect 5499 21502 5555 21511
rect 5931 21567 5987 21576
rect 5931 21502 5987 21511
rect 6275 21555 6331 21564
rect 6275 21490 6331 21499
rect 6699 21555 6755 21564
rect 6699 21490 6755 21499
rect 6275 21161 6331 21170
rect 5027 21149 5083 21158
rect 5027 21084 5083 21093
rect 5499 21149 5555 21158
rect 5499 21084 5555 21093
rect 5931 21149 5987 21158
rect 6275 21096 6331 21105
rect 6699 21161 6755 21170
rect 6699 21096 6755 21105
rect 5931 21084 5987 21093
rect 5027 20777 5083 20786
rect 5027 20712 5083 20721
rect 5499 20777 5555 20786
rect 5499 20712 5555 20721
rect 5931 20777 5987 20786
rect 5931 20712 5987 20721
rect 6275 20765 6331 20774
rect 6275 20700 6331 20709
rect 6699 20765 6755 20774
rect 6699 20700 6755 20709
rect 6275 20371 6331 20380
rect 5027 20359 5083 20368
rect 5027 20294 5083 20303
rect 5499 20359 5555 20368
rect 5499 20294 5555 20303
rect 5931 20359 5987 20368
rect 6275 20306 6331 20315
rect 6699 20371 6755 20380
rect 6699 20306 6755 20315
rect 5931 20294 5987 20303
rect 5027 19987 5083 19996
rect 5027 19922 5083 19931
rect 5499 19987 5555 19996
rect 5499 19922 5555 19931
rect 5931 19987 5987 19996
rect 5931 19922 5987 19931
rect 6275 19975 6331 19984
rect 6275 19910 6331 19919
rect 6699 19975 6755 19984
rect 6699 19910 6755 19919
rect 6275 19581 6331 19590
rect 5027 19569 5083 19578
rect 5027 19504 5083 19513
rect 5499 19569 5555 19578
rect 5499 19504 5555 19513
rect 5931 19569 5987 19578
rect 6275 19516 6331 19525
rect 6699 19581 6755 19590
rect 6699 19516 6755 19525
rect 5931 19504 5987 19513
rect 5027 19197 5083 19206
rect 5027 19132 5083 19141
rect 5499 19197 5555 19206
rect 5499 19132 5555 19141
rect 5931 19197 5987 19206
rect 5931 19132 5987 19141
rect 6275 19185 6331 19194
rect 6275 19120 6331 19129
rect 6699 19185 6755 19194
rect 6699 19120 6755 19129
rect 6275 18791 6331 18800
rect 5027 18779 5083 18788
rect 5027 18714 5083 18723
rect 5499 18779 5555 18788
rect 5499 18714 5555 18723
rect 5931 18779 5987 18788
rect 6275 18726 6331 18735
rect 6699 18791 6755 18800
rect 6699 18726 6755 18735
rect 5931 18714 5987 18723
rect 5027 18407 5083 18416
rect 5027 18342 5083 18351
rect 5499 18407 5555 18416
rect 5499 18342 5555 18351
rect 5931 18407 5987 18416
rect 5931 18342 5987 18351
rect 6275 18395 6331 18404
rect 6275 18330 6331 18339
rect 6699 18395 6755 18404
rect 6699 18330 6755 18339
rect 6275 18001 6331 18010
rect 5027 17989 5083 17998
rect 5027 17924 5083 17933
rect 5499 17989 5555 17998
rect 5499 17924 5555 17933
rect 5931 17989 5987 17998
rect 6275 17936 6331 17945
rect 6699 18001 6755 18010
rect 6699 17936 6755 17945
rect 5931 17924 5987 17933
rect 5027 17617 5083 17626
rect 5027 17552 5083 17561
rect 5499 17617 5555 17626
rect 5499 17552 5555 17561
rect 5931 17617 5987 17626
rect 5931 17552 5987 17561
rect 6275 17605 6331 17614
rect 6275 17540 6331 17549
rect 6699 17605 6755 17614
rect 6699 17540 6755 17549
rect 6275 17211 6331 17220
rect 5027 17199 5083 17208
rect 5027 17134 5083 17143
rect 5499 17199 5555 17208
rect 5499 17134 5555 17143
rect 5931 17199 5987 17208
rect 6275 17146 6331 17155
rect 6699 17211 6755 17220
rect 6699 17146 6755 17155
rect 5931 17134 5987 17143
rect 5027 16827 5083 16836
rect 5027 16762 5083 16771
rect 5499 16827 5555 16836
rect 5499 16762 5555 16771
rect 5931 16827 5987 16836
rect 5931 16762 5987 16771
rect 6275 16815 6331 16824
rect 6275 16750 6331 16759
rect 6699 16815 6755 16824
rect 6699 16750 6755 16759
rect 6275 16421 6331 16430
rect 5027 16409 5083 16418
rect 5027 16344 5083 16353
rect 5499 16409 5555 16418
rect 5499 16344 5555 16353
rect 5931 16409 5987 16418
rect 6275 16356 6331 16365
rect 6699 16421 6755 16430
rect 6699 16356 6755 16365
rect 5931 16344 5987 16353
rect 5027 16037 5083 16046
rect 5027 15972 5083 15981
rect 5499 16037 5555 16046
rect 5499 15972 5555 15981
rect 5931 16037 5987 16046
rect 5931 15972 5987 15981
rect 6275 16025 6331 16034
rect 6275 15960 6331 15969
rect 6699 16025 6755 16034
rect 6699 15960 6755 15969
rect 6275 15631 6331 15640
rect 5027 15619 5083 15628
rect 5027 15554 5083 15563
rect 5499 15619 5555 15628
rect 5499 15554 5555 15563
rect 5931 15619 5987 15628
rect 6275 15566 6331 15575
rect 6699 15631 6755 15640
rect 6699 15566 6755 15575
rect 5931 15554 5987 15563
rect 5027 15247 5083 15256
rect 5027 15182 5083 15191
rect 5499 15247 5555 15256
rect 5499 15182 5555 15191
rect 5931 15247 5987 15256
rect 5931 15182 5987 15191
rect 6275 15235 6331 15244
rect 6275 15170 6331 15179
rect 6699 15235 6755 15244
rect 6699 15170 6755 15179
rect 6275 14841 6331 14850
rect 5027 14829 5083 14838
rect 5027 14764 5083 14773
rect 5499 14829 5555 14838
rect 5499 14764 5555 14773
rect 5931 14829 5987 14838
rect 6275 14776 6331 14785
rect 6699 14841 6755 14850
rect 6699 14776 6755 14785
rect 5931 14764 5987 14773
rect 5027 14457 5083 14466
rect 5027 14392 5083 14401
rect 5499 14457 5555 14466
rect 5499 14392 5555 14401
rect 5931 14457 5987 14466
rect 5931 14392 5987 14401
rect 6275 14445 6331 14454
rect 6275 14380 6331 14389
rect 6699 14445 6755 14454
rect 6699 14380 6755 14389
rect 6275 14051 6331 14060
rect 5027 14039 5083 14048
rect 5027 13974 5083 13983
rect 5499 14039 5555 14048
rect 5499 13974 5555 13983
rect 5931 14039 5987 14048
rect 6275 13986 6331 13995
rect 6699 14051 6755 14060
rect 6699 13986 6755 13995
rect 5931 13974 5987 13983
rect 5027 13667 5083 13676
rect 5027 13602 5083 13611
rect 5499 13667 5555 13676
rect 5499 13602 5555 13611
rect 5931 13667 5987 13676
rect 5931 13602 5987 13611
rect 6275 13655 6331 13664
rect 6275 13590 6331 13599
rect 6699 13655 6755 13664
rect 6699 13590 6755 13599
rect 6275 13261 6331 13270
rect 5027 13249 5083 13258
rect 5027 13184 5083 13193
rect 5499 13249 5555 13258
rect 5499 13184 5555 13193
rect 5931 13249 5987 13258
rect 6275 13196 6331 13205
rect 6699 13261 6755 13270
rect 6699 13196 6755 13205
rect 5931 13184 5987 13193
rect 5027 12877 5083 12886
rect 5027 12812 5083 12821
rect 5499 12877 5555 12886
rect 5499 12812 5555 12821
rect 5931 12877 5987 12886
rect 5931 12812 5987 12821
rect 6275 12865 6331 12874
rect 6275 12800 6331 12809
rect 6699 12865 6755 12874
rect 6699 12800 6755 12809
rect 6275 12471 6331 12480
rect 5027 12459 5083 12468
rect 5027 12394 5083 12403
rect 5499 12459 5555 12468
rect 5499 12394 5555 12403
rect 5931 12459 5987 12468
rect 6275 12406 6331 12415
rect 6699 12471 6755 12480
rect 6699 12406 6755 12415
rect 5931 12394 5987 12403
rect 5027 12087 5083 12096
rect 5027 12022 5083 12031
rect 5499 12087 5555 12096
rect 5499 12022 5555 12031
rect 5931 12087 5987 12096
rect 5931 12022 5987 12031
rect 6275 12075 6331 12084
rect 6275 12010 6331 12019
rect 6699 12075 6755 12084
rect 6699 12010 6755 12019
rect 6275 11681 6331 11690
rect 5027 11669 5083 11678
rect 5027 11604 5083 11613
rect 5499 11669 5555 11678
rect 5499 11604 5555 11613
rect 5931 11669 5987 11678
rect 6275 11616 6331 11625
rect 6699 11681 6755 11690
rect 6699 11616 6755 11625
rect 5931 11604 5987 11613
rect 5027 11297 5083 11306
rect 5027 11232 5083 11241
rect 5499 11297 5555 11306
rect 5499 11232 5555 11241
rect 5931 11297 5987 11306
rect 5931 11232 5987 11241
rect 6275 11285 6331 11294
rect 6275 11220 6331 11229
rect 6699 11285 6755 11294
rect 6699 11220 6755 11229
rect 6275 10891 6331 10900
rect 5027 10879 5083 10888
rect 5027 10814 5083 10823
rect 5499 10879 5555 10888
rect 5499 10814 5555 10823
rect 5931 10879 5987 10888
rect 6275 10826 6331 10835
rect 6699 10891 6755 10900
rect 6699 10826 6755 10835
rect 5931 10814 5987 10823
rect 5027 10507 5083 10516
rect 5027 10442 5083 10451
rect 5499 10507 5555 10516
rect 5499 10442 5555 10451
rect 5931 10507 5987 10516
rect 5931 10442 5987 10451
rect 6275 10495 6331 10504
rect 6275 10430 6331 10439
rect 6699 10495 6755 10504
rect 6699 10430 6755 10439
rect 6275 10101 6331 10110
rect 5027 10089 5083 10098
rect 5027 10024 5083 10033
rect 5499 10089 5555 10098
rect 5499 10024 5555 10033
rect 5931 10089 5987 10098
rect 6275 10036 6331 10045
rect 6699 10101 6755 10110
rect 6699 10036 6755 10045
rect 5931 10024 5987 10033
rect 5027 9717 5083 9726
rect 5027 9652 5083 9661
rect 5499 9717 5555 9726
rect 5499 9652 5555 9661
rect 5931 9717 5987 9726
rect 5931 9652 5987 9661
rect 6275 9705 6331 9714
rect 6275 9640 6331 9649
rect 6699 9705 6755 9714
rect 6699 9640 6755 9649
rect 6275 9311 6331 9320
rect 5027 9299 5083 9308
rect 5027 9234 5083 9243
rect 5499 9299 5555 9308
rect 5499 9234 5555 9243
rect 5931 9299 5987 9308
rect 6275 9246 6331 9255
rect 6699 9311 6755 9320
rect 6699 9246 6755 9255
rect 5931 9234 5987 9243
rect 5027 8927 5083 8936
rect 5027 8862 5083 8871
rect 5499 8927 5555 8936
rect 5499 8862 5555 8871
rect 5931 8927 5987 8936
rect 5931 8862 5987 8871
rect 6275 8915 6331 8924
rect 6275 8850 6331 8859
rect 6699 8915 6755 8924
rect 6699 8850 6755 8859
rect 6275 8521 6331 8530
rect 5027 8509 5083 8518
rect 5027 8444 5083 8453
rect 5499 8509 5555 8518
rect 5499 8444 5555 8453
rect 5931 8509 5987 8518
rect 6275 8456 6331 8465
rect 6699 8521 6755 8530
rect 6699 8456 6755 8465
rect 5931 8444 5987 8453
rect 5027 8137 5083 8146
rect 5027 8072 5083 8081
rect 5499 8137 5555 8146
rect 5499 8072 5555 8081
rect 5931 8137 5987 8146
rect 5931 8072 5987 8081
rect 6275 8125 6331 8134
rect 6275 8060 6331 8069
rect 6699 8125 6755 8134
rect 6699 8060 6755 8069
rect 6275 7731 6331 7740
rect 5027 7719 5083 7728
rect 5027 7654 5083 7663
rect 5499 7719 5555 7728
rect 5499 7654 5555 7663
rect 5931 7719 5987 7728
rect 6275 7666 6331 7675
rect 6699 7731 6755 7740
rect 6699 7666 6755 7675
rect 5931 7654 5987 7663
rect 5027 7347 5083 7356
rect 5027 7282 5083 7291
rect 5499 7347 5555 7356
rect 5499 7282 5555 7291
rect 5931 7347 5987 7356
rect 5931 7282 5987 7291
rect 6275 7335 6331 7344
rect 6275 7270 6331 7279
rect 6699 7335 6755 7344
rect 6699 7270 6755 7279
rect 6275 6941 6331 6950
rect 5027 6929 5083 6938
rect 5027 6864 5083 6873
rect 5499 6929 5555 6938
rect 5499 6864 5555 6873
rect 5931 6929 5987 6938
rect 6275 6876 6331 6885
rect 6699 6941 6755 6950
rect 6699 6876 6755 6885
rect 5931 6864 5987 6873
rect 5027 6557 5083 6566
rect 5027 6492 5083 6501
rect 5499 6557 5555 6566
rect 5499 6492 5555 6501
rect 5931 6557 5987 6566
rect 5931 6492 5987 6501
rect 6275 6545 6331 6554
rect 6275 6480 6331 6489
rect 6699 6545 6755 6554
rect 6699 6480 6755 6489
rect 3661 6226 3713 6232
rect 3661 6168 3713 6174
rect 3673 5939 3701 6168
rect 6275 6151 6331 6160
rect 5027 6139 5083 6148
rect 5027 6074 5083 6083
rect 5499 6139 5555 6148
rect 5499 6074 5555 6083
rect 5931 6139 5987 6148
rect 6275 6086 6331 6095
rect 6699 6151 6755 6160
rect 6699 6086 6755 6095
rect 5931 6074 5987 6083
rect 4629 5939 4635 5951
rect 3673 5911 4635 5939
rect 4629 5899 4635 5911
rect 4687 5899 4693 5951
rect 5027 5767 5083 5776
rect 5027 5702 5083 5711
rect 5499 5767 5555 5776
rect 5499 5702 5555 5711
rect 5931 5767 5987 5776
rect 5931 5702 5987 5711
rect 6275 5755 6331 5764
rect 6275 5690 6331 5699
rect 6699 5755 6755 5764
rect 6699 5690 6755 5699
rect 3661 5676 3713 5682
rect 3661 5618 3713 5624
rect 3673 5544 3701 5618
rect 4549 5544 4555 5556
rect 3673 5516 4555 5544
rect 4549 5504 4555 5516
rect 4607 5504 4613 5556
rect 3661 5436 3713 5442
rect 3661 5378 3713 5384
rect 3673 5149 3701 5378
rect 6275 5361 6331 5370
rect 5027 5349 5083 5358
rect 5027 5284 5083 5293
rect 5499 5349 5555 5358
rect 5499 5284 5555 5293
rect 5931 5349 5987 5358
rect 6275 5296 6331 5305
rect 6699 5361 6755 5370
rect 6699 5296 6755 5305
rect 5931 5284 5987 5293
rect 4469 5149 4475 5161
rect 3673 5121 4475 5149
rect 4469 5109 4475 5121
rect 4527 5109 4533 5161
rect 5027 4977 5083 4986
rect 5027 4912 5083 4921
rect 5499 4977 5555 4986
rect 5499 4912 5555 4921
rect 5931 4977 5987 4986
rect 5931 4912 5987 4921
rect 6275 4965 6331 4974
rect 6275 4900 6331 4909
rect 6699 4965 6755 4974
rect 6699 4900 6755 4909
rect 3661 4886 3713 4892
rect 3661 4828 3713 4834
rect 3673 4754 3701 4828
rect 4389 4754 4395 4766
rect 3673 4726 4395 4754
rect 4389 4714 4395 4726
rect 4447 4714 4453 4766
rect 6275 4571 6331 4580
rect 5027 4559 5083 4568
rect 5027 4494 5083 4503
rect 5499 4559 5555 4568
rect 5499 4494 5555 4503
rect 5931 4559 5987 4568
rect 6275 4506 6331 4515
rect 6699 4571 6755 4580
rect 6699 4506 6755 4515
rect 5931 4494 5987 4503
rect 5027 4187 5083 4196
rect 5027 4122 5083 4131
rect 5499 4187 5555 4196
rect 5499 4122 5555 4131
rect 5931 4187 5987 4196
rect 5931 4122 5987 4131
rect 6275 4175 6331 4184
rect 6275 4110 6331 4119
rect 6699 4175 6755 4184
rect 6699 4110 6755 4119
rect 3661 3856 3713 3862
rect 3661 3798 3713 3804
rect 3673 3569 3701 3798
rect 6275 3781 6331 3790
rect 5027 3769 5083 3778
rect 5027 3704 5083 3713
rect 5499 3769 5555 3778
rect 5499 3704 5555 3713
rect 5931 3769 5987 3778
rect 6275 3716 6331 3725
rect 6699 3781 6755 3790
rect 6699 3716 6755 3725
rect 5931 3704 5987 3713
rect 4309 3569 4315 3581
rect 3673 3541 4315 3569
rect 4309 3529 4315 3541
rect 4367 3529 4373 3581
rect 5027 3397 5083 3406
rect 5027 3332 5083 3341
rect 5499 3397 5555 3406
rect 5499 3332 5555 3341
rect 5931 3397 5987 3406
rect 5931 3332 5987 3341
rect 6275 3385 6331 3394
rect 6275 3320 6331 3329
rect 6699 3385 6755 3394
rect 6699 3320 6755 3329
rect 3661 3306 3713 3312
rect 3661 3248 3713 3254
rect 3673 3174 3701 3248
rect 4229 3174 4235 3186
rect 3673 3146 4235 3174
rect 4229 3134 4235 3146
rect 4287 3134 4293 3186
rect 3661 3066 3713 3072
rect 3661 3008 3713 3014
rect 3673 2779 3701 3008
rect 6275 2991 6331 3000
rect 5027 2979 5083 2988
rect 5027 2914 5083 2923
rect 5499 2979 5555 2988
rect 5499 2914 5555 2923
rect 5931 2979 5987 2988
rect 6275 2926 6331 2935
rect 6699 2991 6755 3000
rect 6699 2926 6755 2935
rect 5931 2914 5987 2923
rect 4149 2779 4155 2791
rect 3673 2751 4155 2779
rect 4149 2739 4155 2751
rect 4207 2739 4213 2791
rect 5027 2607 5083 2616
rect 5027 2542 5083 2551
rect 5499 2607 5555 2616
rect 5499 2542 5555 2551
rect 5931 2607 5987 2616
rect 5931 2542 5987 2551
rect 6275 2595 6331 2604
rect 6275 2530 6331 2539
rect 6699 2595 6755 2604
rect 6699 2530 6755 2539
rect 3661 2516 3713 2522
rect 3661 2458 3713 2464
rect 3673 2384 3701 2458
rect 4069 2384 4075 2396
rect 3673 2356 4075 2384
rect 4069 2344 4075 2356
rect 4127 2344 4133 2396
rect 6275 2201 6331 2210
rect 5027 2189 5083 2198
rect 5027 2124 5083 2133
rect 5499 2189 5555 2198
rect 5499 2124 5555 2133
rect 5931 2189 5987 2198
rect 6275 2136 6331 2145
rect 6699 2201 6755 2210
rect 6699 2136 6755 2145
rect 5931 2124 5987 2133
rect 5027 1817 5083 1826
rect 5027 1752 5083 1761
rect 5499 1817 5555 1826
rect 5499 1752 5555 1761
rect 5931 1817 5987 1826
rect 5931 1752 5987 1761
rect 6275 1805 6331 1814
rect 6275 1740 6331 1749
rect 6699 1805 6755 1814
rect 6699 1740 6755 1749
rect 3661 1486 3713 1492
rect 3661 1428 3713 1434
rect 3673 1199 3701 1428
rect 6275 1411 6331 1420
rect 5027 1399 5083 1408
rect 5027 1334 5083 1343
rect 5499 1399 5555 1408
rect 5499 1334 5555 1343
rect 5931 1399 5987 1408
rect 6275 1346 6331 1355
rect 6699 1411 6755 1420
rect 6699 1346 6755 1355
rect 5931 1334 5987 1343
rect 3989 1199 3995 1211
rect 3673 1171 3995 1199
rect 3989 1159 3995 1171
rect 4047 1159 4053 1211
rect 5027 1027 5083 1036
rect 3909 1013 3915 1025
rect 3673 985 3915 1013
rect 3673 942 3701 985
rect 3909 973 3915 985
rect 3967 973 3973 1025
rect 5027 962 5083 971
rect 5499 1027 5555 1036
rect 5499 962 5555 971
rect 5931 1027 5987 1036
rect 5931 962 5987 971
rect 6275 1015 6331 1024
rect 6275 950 6331 959
rect 6699 1015 6755 1024
rect 6699 950 6755 959
rect 3661 936 3713 942
rect 3661 878 3713 884
rect 3661 696 3713 702
rect 3661 638 3713 644
rect 3673 409 3701 638
rect 6275 621 6331 630
rect 5027 609 5083 618
rect 5027 544 5083 553
rect 5499 609 5555 618
rect 5499 544 5555 553
rect 5931 609 5987 618
rect 6275 556 6331 565
rect 6699 621 6755 630
rect 6699 556 6755 565
rect 5931 544 5987 553
rect 3829 409 3835 421
rect 3673 381 3835 409
rect 3829 369 3835 381
rect 3887 369 3893 421
rect 5027 237 5083 246
rect 3749 223 3755 235
rect 3673 195 3755 223
rect 3673 152 3701 195
rect 3749 183 3755 195
rect 3807 183 3813 235
rect 5027 172 5083 181
rect 5499 237 5555 246
rect 5499 172 5555 181
rect 5931 237 5987 246
rect 5931 172 5987 181
rect 6275 225 6331 234
rect 6275 160 6331 169
rect 6699 225 6755 234
rect 6699 160 6755 169
rect 3661 146 3713 152
rect 3661 88 3713 94
<< via2 >>
rect 6275 25108 6331 25111
rect 5027 25097 5083 25099
rect 5027 25045 5029 25097
rect 5029 25045 5081 25097
rect 5081 25045 5083 25097
rect 5027 25043 5083 25045
rect 5499 25097 5555 25099
rect 5499 25045 5501 25097
rect 5501 25045 5553 25097
rect 5553 25045 5555 25097
rect 5499 25043 5555 25045
rect 5931 25097 5987 25099
rect 5931 25045 5933 25097
rect 5933 25045 5985 25097
rect 5985 25045 5987 25097
rect 6275 25056 6277 25108
rect 6277 25056 6329 25108
rect 6329 25056 6331 25108
rect 6275 25055 6331 25056
rect 6699 25108 6755 25111
rect 6699 25056 6701 25108
rect 6701 25056 6753 25108
rect 6753 25056 6755 25108
rect 6699 25055 6755 25056
rect 5931 25043 5987 25045
rect 5027 24725 5083 24727
rect 5027 24673 5029 24725
rect 5029 24673 5081 24725
rect 5081 24673 5083 24725
rect 5027 24671 5083 24673
rect 5499 24725 5555 24727
rect 5499 24673 5501 24725
rect 5501 24673 5553 24725
rect 5553 24673 5555 24725
rect 5499 24671 5555 24673
rect 5931 24725 5987 24727
rect 5931 24673 5933 24725
rect 5933 24673 5985 24725
rect 5985 24673 5987 24725
rect 5931 24671 5987 24673
rect 6275 24714 6331 24715
rect 6275 24662 6277 24714
rect 6277 24662 6329 24714
rect 6329 24662 6331 24714
rect 6275 24659 6331 24662
rect 6699 24714 6755 24715
rect 6699 24662 6701 24714
rect 6701 24662 6753 24714
rect 6753 24662 6755 24714
rect 6699 24659 6755 24662
rect 6275 24318 6331 24321
rect 5027 24307 5083 24309
rect 5027 24255 5029 24307
rect 5029 24255 5081 24307
rect 5081 24255 5083 24307
rect 5027 24253 5083 24255
rect 5499 24307 5555 24309
rect 5499 24255 5501 24307
rect 5501 24255 5553 24307
rect 5553 24255 5555 24307
rect 5499 24253 5555 24255
rect 5931 24307 5987 24309
rect 5931 24255 5933 24307
rect 5933 24255 5985 24307
rect 5985 24255 5987 24307
rect 6275 24266 6277 24318
rect 6277 24266 6329 24318
rect 6329 24266 6331 24318
rect 6275 24265 6331 24266
rect 6699 24318 6755 24321
rect 6699 24266 6701 24318
rect 6701 24266 6753 24318
rect 6753 24266 6755 24318
rect 6699 24265 6755 24266
rect 5931 24253 5987 24255
rect 5027 23935 5083 23937
rect 5027 23883 5029 23935
rect 5029 23883 5081 23935
rect 5081 23883 5083 23935
rect 5027 23881 5083 23883
rect 5499 23935 5555 23937
rect 5499 23883 5501 23935
rect 5501 23883 5553 23935
rect 5553 23883 5555 23935
rect 5499 23881 5555 23883
rect 5931 23935 5987 23937
rect 5931 23883 5933 23935
rect 5933 23883 5985 23935
rect 5985 23883 5987 23935
rect 5931 23881 5987 23883
rect 6275 23924 6331 23925
rect 6275 23872 6277 23924
rect 6277 23872 6329 23924
rect 6329 23872 6331 23924
rect 6275 23869 6331 23872
rect 6699 23924 6755 23925
rect 6699 23872 6701 23924
rect 6701 23872 6753 23924
rect 6753 23872 6755 23924
rect 6699 23869 6755 23872
rect 6275 23528 6331 23531
rect 5027 23517 5083 23519
rect 5027 23465 5029 23517
rect 5029 23465 5081 23517
rect 5081 23465 5083 23517
rect 5027 23463 5083 23465
rect 5499 23517 5555 23519
rect 5499 23465 5501 23517
rect 5501 23465 5553 23517
rect 5553 23465 5555 23517
rect 5499 23463 5555 23465
rect 5931 23517 5987 23519
rect 5931 23465 5933 23517
rect 5933 23465 5985 23517
rect 5985 23465 5987 23517
rect 6275 23476 6277 23528
rect 6277 23476 6329 23528
rect 6329 23476 6331 23528
rect 6275 23475 6331 23476
rect 6699 23528 6755 23531
rect 6699 23476 6701 23528
rect 6701 23476 6753 23528
rect 6753 23476 6755 23528
rect 6699 23475 6755 23476
rect 5931 23463 5987 23465
rect 5027 23145 5083 23147
rect 5027 23093 5029 23145
rect 5029 23093 5081 23145
rect 5081 23093 5083 23145
rect 5027 23091 5083 23093
rect 5499 23145 5555 23147
rect 5499 23093 5501 23145
rect 5501 23093 5553 23145
rect 5553 23093 5555 23145
rect 5499 23091 5555 23093
rect 5931 23145 5987 23147
rect 5931 23093 5933 23145
rect 5933 23093 5985 23145
rect 5985 23093 5987 23145
rect 5931 23091 5987 23093
rect 6275 23134 6331 23135
rect 6275 23082 6277 23134
rect 6277 23082 6329 23134
rect 6329 23082 6331 23134
rect 6275 23079 6331 23082
rect 6699 23134 6755 23135
rect 6699 23082 6701 23134
rect 6701 23082 6753 23134
rect 6753 23082 6755 23134
rect 6699 23079 6755 23082
rect 6275 22738 6331 22741
rect 5027 22727 5083 22729
rect 5027 22675 5029 22727
rect 5029 22675 5081 22727
rect 5081 22675 5083 22727
rect 5027 22673 5083 22675
rect 5499 22727 5555 22729
rect 5499 22675 5501 22727
rect 5501 22675 5553 22727
rect 5553 22675 5555 22727
rect 5499 22673 5555 22675
rect 5931 22727 5987 22729
rect 5931 22675 5933 22727
rect 5933 22675 5985 22727
rect 5985 22675 5987 22727
rect 6275 22686 6277 22738
rect 6277 22686 6329 22738
rect 6329 22686 6331 22738
rect 6275 22685 6331 22686
rect 6699 22738 6755 22741
rect 6699 22686 6701 22738
rect 6701 22686 6753 22738
rect 6753 22686 6755 22738
rect 6699 22685 6755 22686
rect 5931 22673 5987 22675
rect 5027 22355 5083 22357
rect 5027 22303 5029 22355
rect 5029 22303 5081 22355
rect 5081 22303 5083 22355
rect 5027 22301 5083 22303
rect 5499 22355 5555 22357
rect 5499 22303 5501 22355
rect 5501 22303 5553 22355
rect 5553 22303 5555 22355
rect 5499 22301 5555 22303
rect 5931 22355 5987 22357
rect 5931 22303 5933 22355
rect 5933 22303 5985 22355
rect 5985 22303 5987 22355
rect 5931 22301 5987 22303
rect 6275 22344 6331 22345
rect 6275 22292 6277 22344
rect 6277 22292 6329 22344
rect 6329 22292 6331 22344
rect 6275 22289 6331 22292
rect 6699 22344 6755 22345
rect 6699 22292 6701 22344
rect 6701 22292 6753 22344
rect 6753 22292 6755 22344
rect 6699 22289 6755 22292
rect 6275 21948 6331 21951
rect 5027 21937 5083 21939
rect 5027 21885 5029 21937
rect 5029 21885 5081 21937
rect 5081 21885 5083 21937
rect 5027 21883 5083 21885
rect 5499 21937 5555 21939
rect 5499 21885 5501 21937
rect 5501 21885 5553 21937
rect 5553 21885 5555 21937
rect 5499 21883 5555 21885
rect 5931 21937 5987 21939
rect 5931 21885 5933 21937
rect 5933 21885 5985 21937
rect 5985 21885 5987 21937
rect 6275 21896 6277 21948
rect 6277 21896 6329 21948
rect 6329 21896 6331 21948
rect 6275 21895 6331 21896
rect 6699 21948 6755 21951
rect 6699 21896 6701 21948
rect 6701 21896 6753 21948
rect 6753 21896 6755 21948
rect 6699 21895 6755 21896
rect 5931 21883 5987 21885
rect 5027 21565 5083 21567
rect 5027 21513 5029 21565
rect 5029 21513 5081 21565
rect 5081 21513 5083 21565
rect 5027 21511 5083 21513
rect 5499 21565 5555 21567
rect 5499 21513 5501 21565
rect 5501 21513 5553 21565
rect 5553 21513 5555 21565
rect 5499 21511 5555 21513
rect 5931 21565 5987 21567
rect 5931 21513 5933 21565
rect 5933 21513 5985 21565
rect 5985 21513 5987 21565
rect 5931 21511 5987 21513
rect 6275 21554 6331 21555
rect 6275 21502 6277 21554
rect 6277 21502 6329 21554
rect 6329 21502 6331 21554
rect 6275 21499 6331 21502
rect 6699 21554 6755 21555
rect 6699 21502 6701 21554
rect 6701 21502 6753 21554
rect 6753 21502 6755 21554
rect 6699 21499 6755 21502
rect 6275 21158 6331 21161
rect 5027 21147 5083 21149
rect 5027 21095 5029 21147
rect 5029 21095 5081 21147
rect 5081 21095 5083 21147
rect 5027 21093 5083 21095
rect 5499 21147 5555 21149
rect 5499 21095 5501 21147
rect 5501 21095 5553 21147
rect 5553 21095 5555 21147
rect 5499 21093 5555 21095
rect 5931 21147 5987 21149
rect 5931 21095 5933 21147
rect 5933 21095 5985 21147
rect 5985 21095 5987 21147
rect 6275 21106 6277 21158
rect 6277 21106 6329 21158
rect 6329 21106 6331 21158
rect 6275 21105 6331 21106
rect 6699 21158 6755 21161
rect 6699 21106 6701 21158
rect 6701 21106 6753 21158
rect 6753 21106 6755 21158
rect 6699 21105 6755 21106
rect 5931 21093 5987 21095
rect 5027 20775 5083 20777
rect 5027 20723 5029 20775
rect 5029 20723 5081 20775
rect 5081 20723 5083 20775
rect 5027 20721 5083 20723
rect 5499 20775 5555 20777
rect 5499 20723 5501 20775
rect 5501 20723 5553 20775
rect 5553 20723 5555 20775
rect 5499 20721 5555 20723
rect 5931 20775 5987 20777
rect 5931 20723 5933 20775
rect 5933 20723 5985 20775
rect 5985 20723 5987 20775
rect 5931 20721 5987 20723
rect 6275 20764 6331 20765
rect 6275 20712 6277 20764
rect 6277 20712 6329 20764
rect 6329 20712 6331 20764
rect 6275 20709 6331 20712
rect 6699 20764 6755 20765
rect 6699 20712 6701 20764
rect 6701 20712 6753 20764
rect 6753 20712 6755 20764
rect 6699 20709 6755 20712
rect 6275 20368 6331 20371
rect 5027 20357 5083 20359
rect 5027 20305 5029 20357
rect 5029 20305 5081 20357
rect 5081 20305 5083 20357
rect 5027 20303 5083 20305
rect 5499 20357 5555 20359
rect 5499 20305 5501 20357
rect 5501 20305 5553 20357
rect 5553 20305 5555 20357
rect 5499 20303 5555 20305
rect 5931 20357 5987 20359
rect 5931 20305 5933 20357
rect 5933 20305 5985 20357
rect 5985 20305 5987 20357
rect 6275 20316 6277 20368
rect 6277 20316 6329 20368
rect 6329 20316 6331 20368
rect 6275 20315 6331 20316
rect 6699 20368 6755 20371
rect 6699 20316 6701 20368
rect 6701 20316 6753 20368
rect 6753 20316 6755 20368
rect 6699 20315 6755 20316
rect 5931 20303 5987 20305
rect 5027 19985 5083 19987
rect 5027 19933 5029 19985
rect 5029 19933 5081 19985
rect 5081 19933 5083 19985
rect 5027 19931 5083 19933
rect 5499 19985 5555 19987
rect 5499 19933 5501 19985
rect 5501 19933 5553 19985
rect 5553 19933 5555 19985
rect 5499 19931 5555 19933
rect 5931 19985 5987 19987
rect 5931 19933 5933 19985
rect 5933 19933 5985 19985
rect 5985 19933 5987 19985
rect 5931 19931 5987 19933
rect 6275 19974 6331 19975
rect 6275 19922 6277 19974
rect 6277 19922 6329 19974
rect 6329 19922 6331 19974
rect 6275 19919 6331 19922
rect 6699 19974 6755 19975
rect 6699 19922 6701 19974
rect 6701 19922 6753 19974
rect 6753 19922 6755 19974
rect 6699 19919 6755 19922
rect 6275 19578 6331 19581
rect 5027 19567 5083 19569
rect 5027 19515 5029 19567
rect 5029 19515 5081 19567
rect 5081 19515 5083 19567
rect 5027 19513 5083 19515
rect 5499 19567 5555 19569
rect 5499 19515 5501 19567
rect 5501 19515 5553 19567
rect 5553 19515 5555 19567
rect 5499 19513 5555 19515
rect 5931 19567 5987 19569
rect 5931 19515 5933 19567
rect 5933 19515 5985 19567
rect 5985 19515 5987 19567
rect 6275 19526 6277 19578
rect 6277 19526 6329 19578
rect 6329 19526 6331 19578
rect 6275 19525 6331 19526
rect 6699 19578 6755 19581
rect 6699 19526 6701 19578
rect 6701 19526 6753 19578
rect 6753 19526 6755 19578
rect 6699 19525 6755 19526
rect 5931 19513 5987 19515
rect 5027 19195 5083 19197
rect 5027 19143 5029 19195
rect 5029 19143 5081 19195
rect 5081 19143 5083 19195
rect 5027 19141 5083 19143
rect 5499 19195 5555 19197
rect 5499 19143 5501 19195
rect 5501 19143 5553 19195
rect 5553 19143 5555 19195
rect 5499 19141 5555 19143
rect 5931 19195 5987 19197
rect 5931 19143 5933 19195
rect 5933 19143 5985 19195
rect 5985 19143 5987 19195
rect 5931 19141 5987 19143
rect 6275 19184 6331 19185
rect 6275 19132 6277 19184
rect 6277 19132 6329 19184
rect 6329 19132 6331 19184
rect 6275 19129 6331 19132
rect 6699 19184 6755 19185
rect 6699 19132 6701 19184
rect 6701 19132 6753 19184
rect 6753 19132 6755 19184
rect 6699 19129 6755 19132
rect 6275 18788 6331 18791
rect 5027 18777 5083 18779
rect 5027 18725 5029 18777
rect 5029 18725 5081 18777
rect 5081 18725 5083 18777
rect 5027 18723 5083 18725
rect 5499 18777 5555 18779
rect 5499 18725 5501 18777
rect 5501 18725 5553 18777
rect 5553 18725 5555 18777
rect 5499 18723 5555 18725
rect 5931 18777 5987 18779
rect 5931 18725 5933 18777
rect 5933 18725 5985 18777
rect 5985 18725 5987 18777
rect 6275 18736 6277 18788
rect 6277 18736 6329 18788
rect 6329 18736 6331 18788
rect 6275 18735 6331 18736
rect 6699 18788 6755 18791
rect 6699 18736 6701 18788
rect 6701 18736 6753 18788
rect 6753 18736 6755 18788
rect 6699 18735 6755 18736
rect 5931 18723 5987 18725
rect 5027 18405 5083 18407
rect 5027 18353 5029 18405
rect 5029 18353 5081 18405
rect 5081 18353 5083 18405
rect 5027 18351 5083 18353
rect 5499 18405 5555 18407
rect 5499 18353 5501 18405
rect 5501 18353 5553 18405
rect 5553 18353 5555 18405
rect 5499 18351 5555 18353
rect 5931 18405 5987 18407
rect 5931 18353 5933 18405
rect 5933 18353 5985 18405
rect 5985 18353 5987 18405
rect 5931 18351 5987 18353
rect 6275 18394 6331 18395
rect 6275 18342 6277 18394
rect 6277 18342 6329 18394
rect 6329 18342 6331 18394
rect 6275 18339 6331 18342
rect 6699 18394 6755 18395
rect 6699 18342 6701 18394
rect 6701 18342 6753 18394
rect 6753 18342 6755 18394
rect 6699 18339 6755 18342
rect 6275 17998 6331 18001
rect 5027 17987 5083 17989
rect 5027 17935 5029 17987
rect 5029 17935 5081 17987
rect 5081 17935 5083 17987
rect 5027 17933 5083 17935
rect 5499 17987 5555 17989
rect 5499 17935 5501 17987
rect 5501 17935 5553 17987
rect 5553 17935 5555 17987
rect 5499 17933 5555 17935
rect 5931 17987 5987 17989
rect 5931 17935 5933 17987
rect 5933 17935 5985 17987
rect 5985 17935 5987 17987
rect 6275 17946 6277 17998
rect 6277 17946 6329 17998
rect 6329 17946 6331 17998
rect 6275 17945 6331 17946
rect 6699 17998 6755 18001
rect 6699 17946 6701 17998
rect 6701 17946 6753 17998
rect 6753 17946 6755 17998
rect 6699 17945 6755 17946
rect 5931 17933 5987 17935
rect 5027 17615 5083 17617
rect 5027 17563 5029 17615
rect 5029 17563 5081 17615
rect 5081 17563 5083 17615
rect 5027 17561 5083 17563
rect 5499 17615 5555 17617
rect 5499 17563 5501 17615
rect 5501 17563 5553 17615
rect 5553 17563 5555 17615
rect 5499 17561 5555 17563
rect 5931 17615 5987 17617
rect 5931 17563 5933 17615
rect 5933 17563 5985 17615
rect 5985 17563 5987 17615
rect 5931 17561 5987 17563
rect 6275 17604 6331 17605
rect 6275 17552 6277 17604
rect 6277 17552 6329 17604
rect 6329 17552 6331 17604
rect 6275 17549 6331 17552
rect 6699 17604 6755 17605
rect 6699 17552 6701 17604
rect 6701 17552 6753 17604
rect 6753 17552 6755 17604
rect 6699 17549 6755 17552
rect 6275 17208 6331 17211
rect 5027 17197 5083 17199
rect 5027 17145 5029 17197
rect 5029 17145 5081 17197
rect 5081 17145 5083 17197
rect 5027 17143 5083 17145
rect 5499 17197 5555 17199
rect 5499 17145 5501 17197
rect 5501 17145 5553 17197
rect 5553 17145 5555 17197
rect 5499 17143 5555 17145
rect 5931 17197 5987 17199
rect 5931 17145 5933 17197
rect 5933 17145 5985 17197
rect 5985 17145 5987 17197
rect 6275 17156 6277 17208
rect 6277 17156 6329 17208
rect 6329 17156 6331 17208
rect 6275 17155 6331 17156
rect 6699 17208 6755 17211
rect 6699 17156 6701 17208
rect 6701 17156 6753 17208
rect 6753 17156 6755 17208
rect 6699 17155 6755 17156
rect 5931 17143 5987 17145
rect 5027 16825 5083 16827
rect 5027 16773 5029 16825
rect 5029 16773 5081 16825
rect 5081 16773 5083 16825
rect 5027 16771 5083 16773
rect 5499 16825 5555 16827
rect 5499 16773 5501 16825
rect 5501 16773 5553 16825
rect 5553 16773 5555 16825
rect 5499 16771 5555 16773
rect 5931 16825 5987 16827
rect 5931 16773 5933 16825
rect 5933 16773 5985 16825
rect 5985 16773 5987 16825
rect 5931 16771 5987 16773
rect 6275 16814 6331 16815
rect 6275 16762 6277 16814
rect 6277 16762 6329 16814
rect 6329 16762 6331 16814
rect 6275 16759 6331 16762
rect 6699 16814 6755 16815
rect 6699 16762 6701 16814
rect 6701 16762 6753 16814
rect 6753 16762 6755 16814
rect 6699 16759 6755 16762
rect 6275 16418 6331 16421
rect 5027 16407 5083 16409
rect 5027 16355 5029 16407
rect 5029 16355 5081 16407
rect 5081 16355 5083 16407
rect 5027 16353 5083 16355
rect 5499 16407 5555 16409
rect 5499 16355 5501 16407
rect 5501 16355 5553 16407
rect 5553 16355 5555 16407
rect 5499 16353 5555 16355
rect 5931 16407 5987 16409
rect 5931 16355 5933 16407
rect 5933 16355 5985 16407
rect 5985 16355 5987 16407
rect 6275 16366 6277 16418
rect 6277 16366 6329 16418
rect 6329 16366 6331 16418
rect 6275 16365 6331 16366
rect 6699 16418 6755 16421
rect 6699 16366 6701 16418
rect 6701 16366 6753 16418
rect 6753 16366 6755 16418
rect 6699 16365 6755 16366
rect 5931 16353 5987 16355
rect 5027 16035 5083 16037
rect 5027 15983 5029 16035
rect 5029 15983 5081 16035
rect 5081 15983 5083 16035
rect 5027 15981 5083 15983
rect 5499 16035 5555 16037
rect 5499 15983 5501 16035
rect 5501 15983 5553 16035
rect 5553 15983 5555 16035
rect 5499 15981 5555 15983
rect 5931 16035 5987 16037
rect 5931 15983 5933 16035
rect 5933 15983 5985 16035
rect 5985 15983 5987 16035
rect 5931 15981 5987 15983
rect 6275 16024 6331 16025
rect 6275 15972 6277 16024
rect 6277 15972 6329 16024
rect 6329 15972 6331 16024
rect 6275 15969 6331 15972
rect 6699 16024 6755 16025
rect 6699 15972 6701 16024
rect 6701 15972 6753 16024
rect 6753 15972 6755 16024
rect 6699 15969 6755 15972
rect 6275 15628 6331 15631
rect 5027 15617 5083 15619
rect 5027 15565 5029 15617
rect 5029 15565 5081 15617
rect 5081 15565 5083 15617
rect 5027 15563 5083 15565
rect 5499 15617 5555 15619
rect 5499 15565 5501 15617
rect 5501 15565 5553 15617
rect 5553 15565 5555 15617
rect 5499 15563 5555 15565
rect 5931 15617 5987 15619
rect 5931 15565 5933 15617
rect 5933 15565 5985 15617
rect 5985 15565 5987 15617
rect 6275 15576 6277 15628
rect 6277 15576 6329 15628
rect 6329 15576 6331 15628
rect 6275 15575 6331 15576
rect 6699 15628 6755 15631
rect 6699 15576 6701 15628
rect 6701 15576 6753 15628
rect 6753 15576 6755 15628
rect 6699 15575 6755 15576
rect 5931 15563 5987 15565
rect 5027 15245 5083 15247
rect 5027 15193 5029 15245
rect 5029 15193 5081 15245
rect 5081 15193 5083 15245
rect 5027 15191 5083 15193
rect 5499 15245 5555 15247
rect 5499 15193 5501 15245
rect 5501 15193 5553 15245
rect 5553 15193 5555 15245
rect 5499 15191 5555 15193
rect 5931 15245 5987 15247
rect 5931 15193 5933 15245
rect 5933 15193 5985 15245
rect 5985 15193 5987 15245
rect 5931 15191 5987 15193
rect 6275 15234 6331 15235
rect 6275 15182 6277 15234
rect 6277 15182 6329 15234
rect 6329 15182 6331 15234
rect 6275 15179 6331 15182
rect 6699 15234 6755 15235
rect 6699 15182 6701 15234
rect 6701 15182 6753 15234
rect 6753 15182 6755 15234
rect 6699 15179 6755 15182
rect 6275 14838 6331 14841
rect 5027 14827 5083 14829
rect 5027 14775 5029 14827
rect 5029 14775 5081 14827
rect 5081 14775 5083 14827
rect 5027 14773 5083 14775
rect 5499 14827 5555 14829
rect 5499 14775 5501 14827
rect 5501 14775 5553 14827
rect 5553 14775 5555 14827
rect 5499 14773 5555 14775
rect 5931 14827 5987 14829
rect 5931 14775 5933 14827
rect 5933 14775 5985 14827
rect 5985 14775 5987 14827
rect 6275 14786 6277 14838
rect 6277 14786 6329 14838
rect 6329 14786 6331 14838
rect 6275 14785 6331 14786
rect 6699 14838 6755 14841
rect 6699 14786 6701 14838
rect 6701 14786 6753 14838
rect 6753 14786 6755 14838
rect 6699 14785 6755 14786
rect 5931 14773 5987 14775
rect 5027 14455 5083 14457
rect 5027 14403 5029 14455
rect 5029 14403 5081 14455
rect 5081 14403 5083 14455
rect 5027 14401 5083 14403
rect 5499 14455 5555 14457
rect 5499 14403 5501 14455
rect 5501 14403 5553 14455
rect 5553 14403 5555 14455
rect 5499 14401 5555 14403
rect 5931 14455 5987 14457
rect 5931 14403 5933 14455
rect 5933 14403 5985 14455
rect 5985 14403 5987 14455
rect 5931 14401 5987 14403
rect 6275 14444 6331 14445
rect 6275 14392 6277 14444
rect 6277 14392 6329 14444
rect 6329 14392 6331 14444
rect 6275 14389 6331 14392
rect 6699 14444 6755 14445
rect 6699 14392 6701 14444
rect 6701 14392 6753 14444
rect 6753 14392 6755 14444
rect 6699 14389 6755 14392
rect 6275 14048 6331 14051
rect 5027 14037 5083 14039
rect 5027 13985 5029 14037
rect 5029 13985 5081 14037
rect 5081 13985 5083 14037
rect 5027 13983 5083 13985
rect 5499 14037 5555 14039
rect 5499 13985 5501 14037
rect 5501 13985 5553 14037
rect 5553 13985 5555 14037
rect 5499 13983 5555 13985
rect 5931 14037 5987 14039
rect 5931 13985 5933 14037
rect 5933 13985 5985 14037
rect 5985 13985 5987 14037
rect 6275 13996 6277 14048
rect 6277 13996 6329 14048
rect 6329 13996 6331 14048
rect 6275 13995 6331 13996
rect 6699 14048 6755 14051
rect 6699 13996 6701 14048
rect 6701 13996 6753 14048
rect 6753 13996 6755 14048
rect 6699 13995 6755 13996
rect 5931 13983 5987 13985
rect 5027 13665 5083 13667
rect 5027 13613 5029 13665
rect 5029 13613 5081 13665
rect 5081 13613 5083 13665
rect 5027 13611 5083 13613
rect 5499 13665 5555 13667
rect 5499 13613 5501 13665
rect 5501 13613 5553 13665
rect 5553 13613 5555 13665
rect 5499 13611 5555 13613
rect 5931 13665 5987 13667
rect 5931 13613 5933 13665
rect 5933 13613 5985 13665
rect 5985 13613 5987 13665
rect 5931 13611 5987 13613
rect 6275 13654 6331 13655
rect 6275 13602 6277 13654
rect 6277 13602 6329 13654
rect 6329 13602 6331 13654
rect 6275 13599 6331 13602
rect 6699 13654 6755 13655
rect 6699 13602 6701 13654
rect 6701 13602 6753 13654
rect 6753 13602 6755 13654
rect 6699 13599 6755 13602
rect 6275 13258 6331 13261
rect 5027 13247 5083 13249
rect 5027 13195 5029 13247
rect 5029 13195 5081 13247
rect 5081 13195 5083 13247
rect 5027 13193 5083 13195
rect 5499 13247 5555 13249
rect 5499 13195 5501 13247
rect 5501 13195 5553 13247
rect 5553 13195 5555 13247
rect 5499 13193 5555 13195
rect 5931 13247 5987 13249
rect 5931 13195 5933 13247
rect 5933 13195 5985 13247
rect 5985 13195 5987 13247
rect 6275 13206 6277 13258
rect 6277 13206 6329 13258
rect 6329 13206 6331 13258
rect 6275 13205 6331 13206
rect 6699 13258 6755 13261
rect 6699 13206 6701 13258
rect 6701 13206 6753 13258
rect 6753 13206 6755 13258
rect 6699 13205 6755 13206
rect 5931 13193 5987 13195
rect 5027 12875 5083 12877
rect 5027 12823 5029 12875
rect 5029 12823 5081 12875
rect 5081 12823 5083 12875
rect 5027 12821 5083 12823
rect 5499 12875 5555 12877
rect 5499 12823 5501 12875
rect 5501 12823 5553 12875
rect 5553 12823 5555 12875
rect 5499 12821 5555 12823
rect 5931 12875 5987 12877
rect 5931 12823 5933 12875
rect 5933 12823 5985 12875
rect 5985 12823 5987 12875
rect 5931 12821 5987 12823
rect 6275 12864 6331 12865
rect 6275 12812 6277 12864
rect 6277 12812 6329 12864
rect 6329 12812 6331 12864
rect 6275 12809 6331 12812
rect 6699 12864 6755 12865
rect 6699 12812 6701 12864
rect 6701 12812 6753 12864
rect 6753 12812 6755 12864
rect 6699 12809 6755 12812
rect 6275 12468 6331 12471
rect 5027 12457 5083 12459
rect 5027 12405 5029 12457
rect 5029 12405 5081 12457
rect 5081 12405 5083 12457
rect 5027 12403 5083 12405
rect 5499 12457 5555 12459
rect 5499 12405 5501 12457
rect 5501 12405 5553 12457
rect 5553 12405 5555 12457
rect 5499 12403 5555 12405
rect 5931 12457 5987 12459
rect 5931 12405 5933 12457
rect 5933 12405 5985 12457
rect 5985 12405 5987 12457
rect 6275 12416 6277 12468
rect 6277 12416 6329 12468
rect 6329 12416 6331 12468
rect 6275 12415 6331 12416
rect 6699 12468 6755 12471
rect 6699 12416 6701 12468
rect 6701 12416 6753 12468
rect 6753 12416 6755 12468
rect 6699 12415 6755 12416
rect 5931 12403 5987 12405
rect 5027 12085 5083 12087
rect 5027 12033 5029 12085
rect 5029 12033 5081 12085
rect 5081 12033 5083 12085
rect 5027 12031 5083 12033
rect 5499 12085 5555 12087
rect 5499 12033 5501 12085
rect 5501 12033 5553 12085
rect 5553 12033 5555 12085
rect 5499 12031 5555 12033
rect 5931 12085 5987 12087
rect 5931 12033 5933 12085
rect 5933 12033 5985 12085
rect 5985 12033 5987 12085
rect 5931 12031 5987 12033
rect 6275 12074 6331 12075
rect 6275 12022 6277 12074
rect 6277 12022 6329 12074
rect 6329 12022 6331 12074
rect 6275 12019 6331 12022
rect 6699 12074 6755 12075
rect 6699 12022 6701 12074
rect 6701 12022 6753 12074
rect 6753 12022 6755 12074
rect 6699 12019 6755 12022
rect 6275 11678 6331 11681
rect 5027 11667 5083 11669
rect 5027 11615 5029 11667
rect 5029 11615 5081 11667
rect 5081 11615 5083 11667
rect 5027 11613 5083 11615
rect 5499 11667 5555 11669
rect 5499 11615 5501 11667
rect 5501 11615 5553 11667
rect 5553 11615 5555 11667
rect 5499 11613 5555 11615
rect 5931 11667 5987 11669
rect 5931 11615 5933 11667
rect 5933 11615 5985 11667
rect 5985 11615 5987 11667
rect 6275 11626 6277 11678
rect 6277 11626 6329 11678
rect 6329 11626 6331 11678
rect 6275 11625 6331 11626
rect 6699 11678 6755 11681
rect 6699 11626 6701 11678
rect 6701 11626 6753 11678
rect 6753 11626 6755 11678
rect 6699 11625 6755 11626
rect 5931 11613 5987 11615
rect 5027 11295 5083 11297
rect 5027 11243 5029 11295
rect 5029 11243 5081 11295
rect 5081 11243 5083 11295
rect 5027 11241 5083 11243
rect 5499 11295 5555 11297
rect 5499 11243 5501 11295
rect 5501 11243 5553 11295
rect 5553 11243 5555 11295
rect 5499 11241 5555 11243
rect 5931 11295 5987 11297
rect 5931 11243 5933 11295
rect 5933 11243 5985 11295
rect 5985 11243 5987 11295
rect 5931 11241 5987 11243
rect 6275 11284 6331 11285
rect 6275 11232 6277 11284
rect 6277 11232 6329 11284
rect 6329 11232 6331 11284
rect 6275 11229 6331 11232
rect 6699 11284 6755 11285
rect 6699 11232 6701 11284
rect 6701 11232 6753 11284
rect 6753 11232 6755 11284
rect 6699 11229 6755 11232
rect 6275 10888 6331 10891
rect 5027 10877 5083 10879
rect 5027 10825 5029 10877
rect 5029 10825 5081 10877
rect 5081 10825 5083 10877
rect 5027 10823 5083 10825
rect 5499 10877 5555 10879
rect 5499 10825 5501 10877
rect 5501 10825 5553 10877
rect 5553 10825 5555 10877
rect 5499 10823 5555 10825
rect 5931 10877 5987 10879
rect 5931 10825 5933 10877
rect 5933 10825 5985 10877
rect 5985 10825 5987 10877
rect 6275 10836 6277 10888
rect 6277 10836 6329 10888
rect 6329 10836 6331 10888
rect 6275 10835 6331 10836
rect 6699 10888 6755 10891
rect 6699 10836 6701 10888
rect 6701 10836 6753 10888
rect 6753 10836 6755 10888
rect 6699 10835 6755 10836
rect 5931 10823 5987 10825
rect 5027 10505 5083 10507
rect 5027 10453 5029 10505
rect 5029 10453 5081 10505
rect 5081 10453 5083 10505
rect 5027 10451 5083 10453
rect 5499 10505 5555 10507
rect 5499 10453 5501 10505
rect 5501 10453 5553 10505
rect 5553 10453 5555 10505
rect 5499 10451 5555 10453
rect 5931 10505 5987 10507
rect 5931 10453 5933 10505
rect 5933 10453 5985 10505
rect 5985 10453 5987 10505
rect 5931 10451 5987 10453
rect 6275 10494 6331 10495
rect 6275 10442 6277 10494
rect 6277 10442 6329 10494
rect 6329 10442 6331 10494
rect 6275 10439 6331 10442
rect 6699 10494 6755 10495
rect 6699 10442 6701 10494
rect 6701 10442 6753 10494
rect 6753 10442 6755 10494
rect 6699 10439 6755 10442
rect 6275 10098 6331 10101
rect 5027 10087 5083 10089
rect 5027 10035 5029 10087
rect 5029 10035 5081 10087
rect 5081 10035 5083 10087
rect 5027 10033 5083 10035
rect 5499 10087 5555 10089
rect 5499 10035 5501 10087
rect 5501 10035 5553 10087
rect 5553 10035 5555 10087
rect 5499 10033 5555 10035
rect 5931 10087 5987 10089
rect 5931 10035 5933 10087
rect 5933 10035 5985 10087
rect 5985 10035 5987 10087
rect 6275 10046 6277 10098
rect 6277 10046 6329 10098
rect 6329 10046 6331 10098
rect 6275 10045 6331 10046
rect 6699 10098 6755 10101
rect 6699 10046 6701 10098
rect 6701 10046 6753 10098
rect 6753 10046 6755 10098
rect 6699 10045 6755 10046
rect 5931 10033 5987 10035
rect 5027 9715 5083 9717
rect 5027 9663 5029 9715
rect 5029 9663 5081 9715
rect 5081 9663 5083 9715
rect 5027 9661 5083 9663
rect 5499 9715 5555 9717
rect 5499 9663 5501 9715
rect 5501 9663 5553 9715
rect 5553 9663 5555 9715
rect 5499 9661 5555 9663
rect 5931 9715 5987 9717
rect 5931 9663 5933 9715
rect 5933 9663 5985 9715
rect 5985 9663 5987 9715
rect 5931 9661 5987 9663
rect 6275 9704 6331 9705
rect 6275 9652 6277 9704
rect 6277 9652 6329 9704
rect 6329 9652 6331 9704
rect 6275 9649 6331 9652
rect 6699 9704 6755 9705
rect 6699 9652 6701 9704
rect 6701 9652 6753 9704
rect 6753 9652 6755 9704
rect 6699 9649 6755 9652
rect 6275 9308 6331 9311
rect 5027 9297 5083 9299
rect 5027 9245 5029 9297
rect 5029 9245 5081 9297
rect 5081 9245 5083 9297
rect 5027 9243 5083 9245
rect 5499 9297 5555 9299
rect 5499 9245 5501 9297
rect 5501 9245 5553 9297
rect 5553 9245 5555 9297
rect 5499 9243 5555 9245
rect 5931 9297 5987 9299
rect 5931 9245 5933 9297
rect 5933 9245 5985 9297
rect 5985 9245 5987 9297
rect 6275 9256 6277 9308
rect 6277 9256 6329 9308
rect 6329 9256 6331 9308
rect 6275 9255 6331 9256
rect 6699 9308 6755 9311
rect 6699 9256 6701 9308
rect 6701 9256 6753 9308
rect 6753 9256 6755 9308
rect 6699 9255 6755 9256
rect 5931 9243 5987 9245
rect 5027 8925 5083 8927
rect 5027 8873 5029 8925
rect 5029 8873 5081 8925
rect 5081 8873 5083 8925
rect 5027 8871 5083 8873
rect 5499 8925 5555 8927
rect 5499 8873 5501 8925
rect 5501 8873 5553 8925
rect 5553 8873 5555 8925
rect 5499 8871 5555 8873
rect 5931 8925 5987 8927
rect 5931 8873 5933 8925
rect 5933 8873 5985 8925
rect 5985 8873 5987 8925
rect 5931 8871 5987 8873
rect 6275 8914 6331 8915
rect 6275 8862 6277 8914
rect 6277 8862 6329 8914
rect 6329 8862 6331 8914
rect 6275 8859 6331 8862
rect 6699 8914 6755 8915
rect 6699 8862 6701 8914
rect 6701 8862 6753 8914
rect 6753 8862 6755 8914
rect 6699 8859 6755 8862
rect 6275 8518 6331 8521
rect 5027 8507 5083 8509
rect 5027 8455 5029 8507
rect 5029 8455 5081 8507
rect 5081 8455 5083 8507
rect 5027 8453 5083 8455
rect 5499 8507 5555 8509
rect 5499 8455 5501 8507
rect 5501 8455 5553 8507
rect 5553 8455 5555 8507
rect 5499 8453 5555 8455
rect 5931 8507 5987 8509
rect 5931 8455 5933 8507
rect 5933 8455 5985 8507
rect 5985 8455 5987 8507
rect 6275 8466 6277 8518
rect 6277 8466 6329 8518
rect 6329 8466 6331 8518
rect 6275 8465 6331 8466
rect 6699 8518 6755 8521
rect 6699 8466 6701 8518
rect 6701 8466 6753 8518
rect 6753 8466 6755 8518
rect 6699 8465 6755 8466
rect 5931 8453 5987 8455
rect 5027 8135 5083 8137
rect 5027 8083 5029 8135
rect 5029 8083 5081 8135
rect 5081 8083 5083 8135
rect 5027 8081 5083 8083
rect 5499 8135 5555 8137
rect 5499 8083 5501 8135
rect 5501 8083 5553 8135
rect 5553 8083 5555 8135
rect 5499 8081 5555 8083
rect 5931 8135 5987 8137
rect 5931 8083 5933 8135
rect 5933 8083 5985 8135
rect 5985 8083 5987 8135
rect 5931 8081 5987 8083
rect 6275 8124 6331 8125
rect 6275 8072 6277 8124
rect 6277 8072 6329 8124
rect 6329 8072 6331 8124
rect 6275 8069 6331 8072
rect 6699 8124 6755 8125
rect 6699 8072 6701 8124
rect 6701 8072 6753 8124
rect 6753 8072 6755 8124
rect 6699 8069 6755 8072
rect 6275 7728 6331 7731
rect 5027 7717 5083 7719
rect 5027 7665 5029 7717
rect 5029 7665 5081 7717
rect 5081 7665 5083 7717
rect 5027 7663 5083 7665
rect 5499 7717 5555 7719
rect 5499 7665 5501 7717
rect 5501 7665 5553 7717
rect 5553 7665 5555 7717
rect 5499 7663 5555 7665
rect 5931 7717 5987 7719
rect 5931 7665 5933 7717
rect 5933 7665 5985 7717
rect 5985 7665 5987 7717
rect 6275 7676 6277 7728
rect 6277 7676 6329 7728
rect 6329 7676 6331 7728
rect 6275 7675 6331 7676
rect 6699 7728 6755 7731
rect 6699 7676 6701 7728
rect 6701 7676 6753 7728
rect 6753 7676 6755 7728
rect 6699 7675 6755 7676
rect 5931 7663 5987 7665
rect 5027 7345 5083 7347
rect 5027 7293 5029 7345
rect 5029 7293 5081 7345
rect 5081 7293 5083 7345
rect 5027 7291 5083 7293
rect 5499 7345 5555 7347
rect 5499 7293 5501 7345
rect 5501 7293 5553 7345
rect 5553 7293 5555 7345
rect 5499 7291 5555 7293
rect 5931 7345 5987 7347
rect 5931 7293 5933 7345
rect 5933 7293 5985 7345
rect 5985 7293 5987 7345
rect 5931 7291 5987 7293
rect 6275 7334 6331 7335
rect 6275 7282 6277 7334
rect 6277 7282 6329 7334
rect 6329 7282 6331 7334
rect 6275 7279 6331 7282
rect 6699 7334 6755 7335
rect 6699 7282 6701 7334
rect 6701 7282 6753 7334
rect 6753 7282 6755 7334
rect 6699 7279 6755 7282
rect 6275 6938 6331 6941
rect 5027 6927 5083 6929
rect 5027 6875 5029 6927
rect 5029 6875 5081 6927
rect 5081 6875 5083 6927
rect 5027 6873 5083 6875
rect 5499 6927 5555 6929
rect 5499 6875 5501 6927
rect 5501 6875 5553 6927
rect 5553 6875 5555 6927
rect 5499 6873 5555 6875
rect 5931 6927 5987 6929
rect 5931 6875 5933 6927
rect 5933 6875 5985 6927
rect 5985 6875 5987 6927
rect 6275 6886 6277 6938
rect 6277 6886 6329 6938
rect 6329 6886 6331 6938
rect 6275 6885 6331 6886
rect 6699 6938 6755 6941
rect 6699 6886 6701 6938
rect 6701 6886 6753 6938
rect 6753 6886 6755 6938
rect 6699 6885 6755 6886
rect 5931 6873 5987 6875
rect 5027 6555 5083 6557
rect 5027 6503 5029 6555
rect 5029 6503 5081 6555
rect 5081 6503 5083 6555
rect 5027 6501 5083 6503
rect 5499 6555 5555 6557
rect 5499 6503 5501 6555
rect 5501 6503 5553 6555
rect 5553 6503 5555 6555
rect 5499 6501 5555 6503
rect 5931 6555 5987 6557
rect 5931 6503 5933 6555
rect 5933 6503 5985 6555
rect 5985 6503 5987 6555
rect 5931 6501 5987 6503
rect 6275 6544 6331 6545
rect 6275 6492 6277 6544
rect 6277 6492 6329 6544
rect 6329 6492 6331 6544
rect 6275 6489 6331 6492
rect 6699 6544 6755 6545
rect 6699 6492 6701 6544
rect 6701 6492 6753 6544
rect 6753 6492 6755 6544
rect 6699 6489 6755 6492
rect 6275 6148 6331 6151
rect 5027 6137 5083 6139
rect 5027 6085 5029 6137
rect 5029 6085 5081 6137
rect 5081 6085 5083 6137
rect 5027 6083 5083 6085
rect 5499 6137 5555 6139
rect 5499 6085 5501 6137
rect 5501 6085 5553 6137
rect 5553 6085 5555 6137
rect 5499 6083 5555 6085
rect 5931 6137 5987 6139
rect 5931 6085 5933 6137
rect 5933 6085 5985 6137
rect 5985 6085 5987 6137
rect 6275 6096 6277 6148
rect 6277 6096 6329 6148
rect 6329 6096 6331 6148
rect 6275 6095 6331 6096
rect 6699 6148 6755 6151
rect 6699 6096 6701 6148
rect 6701 6096 6753 6148
rect 6753 6096 6755 6148
rect 6699 6095 6755 6096
rect 5931 6083 5987 6085
rect 5027 5765 5083 5767
rect 5027 5713 5029 5765
rect 5029 5713 5081 5765
rect 5081 5713 5083 5765
rect 5027 5711 5083 5713
rect 5499 5765 5555 5767
rect 5499 5713 5501 5765
rect 5501 5713 5553 5765
rect 5553 5713 5555 5765
rect 5499 5711 5555 5713
rect 5931 5765 5987 5767
rect 5931 5713 5933 5765
rect 5933 5713 5985 5765
rect 5985 5713 5987 5765
rect 5931 5711 5987 5713
rect 6275 5754 6331 5755
rect 6275 5702 6277 5754
rect 6277 5702 6329 5754
rect 6329 5702 6331 5754
rect 6275 5699 6331 5702
rect 6699 5754 6755 5755
rect 6699 5702 6701 5754
rect 6701 5702 6753 5754
rect 6753 5702 6755 5754
rect 6699 5699 6755 5702
rect 6275 5358 6331 5361
rect 5027 5347 5083 5349
rect 5027 5295 5029 5347
rect 5029 5295 5081 5347
rect 5081 5295 5083 5347
rect 5027 5293 5083 5295
rect 5499 5347 5555 5349
rect 5499 5295 5501 5347
rect 5501 5295 5553 5347
rect 5553 5295 5555 5347
rect 5499 5293 5555 5295
rect 5931 5347 5987 5349
rect 5931 5295 5933 5347
rect 5933 5295 5985 5347
rect 5985 5295 5987 5347
rect 6275 5306 6277 5358
rect 6277 5306 6329 5358
rect 6329 5306 6331 5358
rect 6275 5305 6331 5306
rect 6699 5358 6755 5361
rect 6699 5306 6701 5358
rect 6701 5306 6753 5358
rect 6753 5306 6755 5358
rect 6699 5305 6755 5306
rect 5931 5293 5987 5295
rect 5027 4975 5083 4977
rect 5027 4923 5029 4975
rect 5029 4923 5081 4975
rect 5081 4923 5083 4975
rect 5027 4921 5083 4923
rect 5499 4975 5555 4977
rect 5499 4923 5501 4975
rect 5501 4923 5553 4975
rect 5553 4923 5555 4975
rect 5499 4921 5555 4923
rect 5931 4975 5987 4977
rect 5931 4923 5933 4975
rect 5933 4923 5985 4975
rect 5985 4923 5987 4975
rect 5931 4921 5987 4923
rect 6275 4964 6331 4965
rect 6275 4912 6277 4964
rect 6277 4912 6329 4964
rect 6329 4912 6331 4964
rect 6275 4909 6331 4912
rect 6699 4964 6755 4965
rect 6699 4912 6701 4964
rect 6701 4912 6753 4964
rect 6753 4912 6755 4964
rect 6699 4909 6755 4912
rect 6275 4568 6331 4571
rect 5027 4557 5083 4559
rect 5027 4505 5029 4557
rect 5029 4505 5081 4557
rect 5081 4505 5083 4557
rect 5027 4503 5083 4505
rect 5499 4557 5555 4559
rect 5499 4505 5501 4557
rect 5501 4505 5553 4557
rect 5553 4505 5555 4557
rect 5499 4503 5555 4505
rect 5931 4557 5987 4559
rect 5931 4505 5933 4557
rect 5933 4505 5985 4557
rect 5985 4505 5987 4557
rect 6275 4516 6277 4568
rect 6277 4516 6329 4568
rect 6329 4516 6331 4568
rect 6275 4515 6331 4516
rect 6699 4568 6755 4571
rect 6699 4516 6701 4568
rect 6701 4516 6753 4568
rect 6753 4516 6755 4568
rect 6699 4515 6755 4516
rect 5931 4503 5987 4505
rect 5027 4185 5083 4187
rect 5027 4133 5029 4185
rect 5029 4133 5081 4185
rect 5081 4133 5083 4185
rect 5027 4131 5083 4133
rect 5499 4185 5555 4187
rect 5499 4133 5501 4185
rect 5501 4133 5553 4185
rect 5553 4133 5555 4185
rect 5499 4131 5555 4133
rect 5931 4185 5987 4187
rect 5931 4133 5933 4185
rect 5933 4133 5985 4185
rect 5985 4133 5987 4185
rect 5931 4131 5987 4133
rect 6275 4174 6331 4175
rect 6275 4122 6277 4174
rect 6277 4122 6329 4174
rect 6329 4122 6331 4174
rect 6275 4119 6331 4122
rect 6699 4174 6755 4175
rect 6699 4122 6701 4174
rect 6701 4122 6753 4174
rect 6753 4122 6755 4174
rect 6699 4119 6755 4122
rect 6275 3778 6331 3781
rect 5027 3767 5083 3769
rect 5027 3715 5029 3767
rect 5029 3715 5081 3767
rect 5081 3715 5083 3767
rect 5027 3713 5083 3715
rect 5499 3767 5555 3769
rect 5499 3715 5501 3767
rect 5501 3715 5553 3767
rect 5553 3715 5555 3767
rect 5499 3713 5555 3715
rect 5931 3767 5987 3769
rect 5931 3715 5933 3767
rect 5933 3715 5985 3767
rect 5985 3715 5987 3767
rect 6275 3726 6277 3778
rect 6277 3726 6329 3778
rect 6329 3726 6331 3778
rect 6275 3725 6331 3726
rect 6699 3778 6755 3781
rect 6699 3726 6701 3778
rect 6701 3726 6753 3778
rect 6753 3726 6755 3778
rect 6699 3725 6755 3726
rect 5931 3713 5987 3715
rect 5027 3395 5083 3397
rect 5027 3343 5029 3395
rect 5029 3343 5081 3395
rect 5081 3343 5083 3395
rect 5027 3341 5083 3343
rect 5499 3395 5555 3397
rect 5499 3343 5501 3395
rect 5501 3343 5553 3395
rect 5553 3343 5555 3395
rect 5499 3341 5555 3343
rect 5931 3395 5987 3397
rect 5931 3343 5933 3395
rect 5933 3343 5985 3395
rect 5985 3343 5987 3395
rect 5931 3341 5987 3343
rect 6275 3384 6331 3385
rect 6275 3332 6277 3384
rect 6277 3332 6329 3384
rect 6329 3332 6331 3384
rect 6275 3329 6331 3332
rect 6699 3384 6755 3385
rect 6699 3332 6701 3384
rect 6701 3332 6753 3384
rect 6753 3332 6755 3384
rect 6699 3329 6755 3332
rect 6275 2988 6331 2991
rect 5027 2977 5083 2979
rect 5027 2925 5029 2977
rect 5029 2925 5081 2977
rect 5081 2925 5083 2977
rect 5027 2923 5083 2925
rect 5499 2977 5555 2979
rect 5499 2925 5501 2977
rect 5501 2925 5553 2977
rect 5553 2925 5555 2977
rect 5499 2923 5555 2925
rect 5931 2977 5987 2979
rect 5931 2925 5933 2977
rect 5933 2925 5985 2977
rect 5985 2925 5987 2977
rect 6275 2936 6277 2988
rect 6277 2936 6329 2988
rect 6329 2936 6331 2988
rect 6275 2935 6331 2936
rect 6699 2988 6755 2991
rect 6699 2936 6701 2988
rect 6701 2936 6753 2988
rect 6753 2936 6755 2988
rect 6699 2935 6755 2936
rect 5931 2923 5987 2925
rect 5027 2605 5083 2607
rect 5027 2553 5029 2605
rect 5029 2553 5081 2605
rect 5081 2553 5083 2605
rect 5027 2551 5083 2553
rect 5499 2605 5555 2607
rect 5499 2553 5501 2605
rect 5501 2553 5553 2605
rect 5553 2553 5555 2605
rect 5499 2551 5555 2553
rect 5931 2605 5987 2607
rect 5931 2553 5933 2605
rect 5933 2553 5985 2605
rect 5985 2553 5987 2605
rect 5931 2551 5987 2553
rect 6275 2594 6331 2595
rect 6275 2542 6277 2594
rect 6277 2542 6329 2594
rect 6329 2542 6331 2594
rect 6275 2539 6331 2542
rect 6699 2594 6755 2595
rect 6699 2542 6701 2594
rect 6701 2542 6753 2594
rect 6753 2542 6755 2594
rect 6699 2539 6755 2542
rect 6275 2198 6331 2201
rect 5027 2187 5083 2189
rect 5027 2135 5029 2187
rect 5029 2135 5081 2187
rect 5081 2135 5083 2187
rect 5027 2133 5083 2135
rect 5499 2187 5555 2189
rect 5499 2135 5501 2187
rect 5501 2135 5553 2187
rect 5553 2135 5555 2187
rect 5499 2133 5555 2135
rect 5931 2187 5987 2189
rect 5931 2135 5933 2187
rect 5933 2135 5985 2187
rect 5985 2135 5987 2187
rect 6275 2146 6277 2198
rect 6277 2146 6329 2198
rect 6329 2146 6331 2198
rect 6275 2145 6331 2146
rect 6699 2198 6755 2201
rect 6699 2146 6701 2198
rect 6701 2146 6753 2198
rect 6753 2146 6755 2198
rect 6699 2145 6755 2146
rect 5931 2133 5987 2135
rect 5027 1815 5083 1817
rect 5027 1763 5029 1815
rect 5029 1763 5081 1815
rect 5081 1763 5083 1815
rect 5027 1761 5083 1763
rect 5499 1815 5555 1817
rect 5499 1763 5501 1815
rect 5501 1763 5553 1815
rect 5553 1763 5555 1815
rect 5499 1761 5555 1763
rect 5931 1815 5987 1817
rect 5931 1763 5933 1815
rect 5933 1763 5985 1815
rect 5985 1763 5987 1815
rect 5931 1761 5987 1763
rect 6275 1804 6331 1805
rect 6275 1752 6277 1804
rect 6277 1752 6329 1804
rect 6329 1752 6331 1804
rect 6275 1749 6331 1752
rect 6699 1804 6755 1805
rect 6699 1752 6701 1804
rect 6701 1752 6753 1804
rect 6753 1752 6755 1804
rect 6699 1749 6755 1752
rect 6275 1408 6331 1411
rect 5027 1397 5083 1399
rect 5027 1345 5029 1397
rect 5029 1345 5081 1397
rect 5081 1345 5083 1397
rect 5027 1343 5083 1345
rect 5499 1397 5555 1399
rect 5499 1345 5501 1397
rect 5501 1345 5553 1397
rect 5553 1345 5555 1397
rect 5499 1343 5555 1345
rect 5931 1397 5987 1399
rect 5931 1345 5933 1397
rect 5933 1345 5985 1397
rect 5985 1345 5987 1397
rect 6275 1356 6277 1408
rect 6277 1356 6329 1408
rect 6329 1356 6331 1408
rect 6275 1355 6331 1356
rect 6699 1408 6755 1411
rect 6699 1356 6701 1408
rect 6701 1356 6753 1408
rect 6753 1356 6755 1408
rect 6699 1355 6755 1356
rect 5931 1343 5987 1345
rect 5027 1025 5083 1027
rect 5027 973 5029 1025
rect 5029 973 5081 1025
rect 5081 973 5083 1025
rect 5027 971 5083 973
rect 5499 1025 5555 1027
rect 5499 973 5501 1025
rect 5501 973 5553 1025
rect 5553 973 5555 1025
rect 5499 971 5555 973
rect 5931 1025 5987 1027
rect 5931 973 5933 1025
rect 5933 973 5985 1025
rect 5985 973 5987 1025
rect 5931 971 5987 973
rect 6275 1014 6331 1015
rect 6275 962 6277 1014
rect 6277 962 6329 1014
rect 6329 962 6331 1014
rect 6275 959 6331 962
rect 6699 1014 6755 1015
rect 6699 962 6701 1014
rect 6701 962 6753 1014
rect 6753 962 6755 1014
rect 6699 959 6755 962
rect 6275 618 6331 621
rect 5027 607 5083 609
rect 5027 555 5029 607
rect 5029 555 5081 607
rect 5081 555 5083 607
rect 5027 553 5083 555
rect 5499 607 5555 609
rect 5499 555 5501 607
rect 5501 555 5553 607
rect 5553 555 5555 607
rect 5499 553 5555 555
rect 5931 607 5987 609
rect 5931 555 5933 607
rect 5933 555 5985 607
rect 5985 555 5987 607
rect 6275 566 6277 618
rect 6277 566 6329 618
rect 6329 566 6331 618
rect 6275 565 6331 566
rect 6699 618 6755 621
rect 6699 566 6701 618
rect 6701 566 6753 618
rect 6753 566 6755 618
rect 6699 565 6755 566
rect 5931 553 5987 555
rect 5027 235 5083 237
rect 5027 183 5029 235
rect 5029 183 5081 235
rect 5081 183 5083 235
rect 5027 181 5083 183
rect 5499 235 5555 237
rect 5499 183 5501 235
rect 5501 183 5553 235
rect 5553 183 5555 235
rect 5499 181 5555 183
rect 5931 235 5987 237
rect 5931 183 5933 235
rect 5933 183 5985 235
rect 5985 183 5987 235
rect 5931 181 5987 183
rect 6275 224 6331 225
rect 6275 172 6277 224
rect 6277 172 6329 224
rect 6329 172 6331 224
rect 6275 169 6331 172
rect 6699 224 6755 225
rect 6699 172 6701 224
rect 6701 172 6753 224
rect 6753 172 6755 224
rect 6699 169 6755 172
<< metal3 >>
rect 6270 25115 6336 25116
rect 6694 25115 6760 25116
rect 6265 25114 6271 25115
rect 5022 25103 5088 25104
rect 5494 25103 5560 25104
rect 5926 25103 5992 25104
rect 4980 25039 5023 25103
rect 5087 25039 5130 25103
rect 5452 25039 5495 25103
rect 5559 25039 5602 25103
rect 5884 25039 5927 25103
rect 5991 25039 6034 25103
rect 6228 25051 6271 25114
rect 6335 25114 6341 25115
rect 6689 25114 6695 25115
rect 6335 25051 6378 25114
rect 6228 25050 6378 25051
rect 6652 25051 6695 25114
rect 6759 25114 6765 25115
rect 6759 25051 6802 25114
rect 6652 25050 6802 25051
rect 5022 25038 5088 25039
rect 5494 25038 5560 25039
rect 5926 25038 5992 25039
rect 5022 24731 5088 24732
rect 5494 24731 5560 24732
rect 5926 24731 5992 24732
rect 4980 24667 5023 24731
rect 5087 24667 5130 24731
rect 5452 24667 5495 24731
rect 5559 24667 5602 24731
rect 5884 24667 5927 24731
rect 5991 24667 6034 24731
rect 6228 24719 6378 24720
rect 5022 24666 5088 24667
rect 5494 24666 5560 24667
rect 5926 24666 5992 24667
rect 6228 24656 6271 24719
rect 6265 24655 6271 24656
rect 6335 24656 6378 24719
rect 6652 24719 6802 24720
rect 6652 24656 6695 24719
rect 6335 24655 6341 24656
rect 6689 24655 6695 24656
rect 6759 24656 6802 24719
rect 6759 24655 6765 24656
rect 6270 24654 6336 24655
rect 6694 24654 6760 24655
rect 6270 24325 6336 24326
rect 6694 24325 6760 24326
rect 6265 24324 6271 24325
rect 5022 24313 5088 24314
rect 5494 24313 5560 24314
rect 5926 24313 5992 24314
rect 4980 24249 5023 24313
rect 5087 24249 5130 24313
rect 5452 24249 5495 24313
rect 5559 24249 5602 24313
rect 5884 24249 5927 24313
rect 5991 24249 6034 24313
rect 6228 24261 6271 24324
rect 6335 24324 6341 24325
rect 6689 24324 6695 24325
rect 6335 24261 6378 24324
rect 6228 24260 6378 24261
rect 6652 24261 6695 24324
rect 6759 24324 6765 24325
rect 6759 24261 6802 24324
rect 6652 24260 6802 24261
rect 5022 24248 5088 24249
rect 5494 24248 5560 24249
rect 5926 24248 5992 24249
rect 5022 23941 5088 23942
rect 5494 23941 5560 23942
rect 5926 23941 5992 23942
rect 4980 23877 5023 23941
rect 5087 23877 5130 23941
rect 5452 23877 5495 23941
rect 5559 23877 5602 23941
rect 5884 23877 5927 23941
rect 5991 23877 6034 23941
rect 6228 23929 6378 23930
rect 5022 23876 5088 23877
rect 5494 23876 5560 23877
rect 5926 23876 5992 23877
rect 6228 23866 6271 23929
rect 6265 23865 6271 23866
rect 6335 23866 6378 23929
rect 6652 23929 6802 23930
rect 6652 23866 6695 23929
rect 6335 23865 6341 23866
rect 6689 23865 6695 23866
rect 6759 23866 6802 23929
rect 6759 23865 6765 23866
rect 6270 23864 6336 23865
rect 6694 23864 6760 23865
rect 6270 23535 6336 23536
rect 6694 23535 6760 23536
rect 6265 23534 6271 23535
rect 5022 23523 5088 23524
rect 5494 23523 5560 23524
rect 5926 23523 5992 23524
rect 4980 23459 5023 23523
rect 5087 23459 5130 23523
rect 5452 23459 5495 23523
rect 5559 23459 5602 23523
rect 5884 23459 5927 23523
rect 5991 23459 6034 23523
rect 6228 23471 6271 23534
rect 6335 23534 6341 23535
rect 6689 23534 6695 23535
rect 6335 23471 6378 23534
rect 6228 23470 6378 23471
rect 6652 23471 6695 23534
rect 6759 23534 6765 23535
rect 6759 23471 6802 23534
rect 6652 23470 6802 23471
rect 5022 23458 5088 23459
rect 5494 23458 5560 23459
rect 5926 23458 5992 23459
rect 5022 23151 5088 23152
rect 5494 23151 5560 23152
rect 5926 23151 5992 23152
rect 4980 23087 5023 23151
rect 5087 23087 5130 23151
rect 5452 23087 5495 23151
rect 5559 23087 5602 23151
rect 5884 23087 5927 23151
rect 5991 23087 6034 23151
rect 6228 23139 6378 23140
rect 5022 23086 5088 23087
rect 5494 23086 5560 23087
rect 5926 23086 5992 23087
rect 6228 23076 6271 23139
rect 6265 23075 6271 23076
rect 6335 23076 6378 23139
rect 6652 23139 6802 23140
rect 6652 23076 6695 23139
rect 6335 23075 6341 23076
rect 6689 23075 6695 23076
rect 6759 23076 6802 23139
rect 6759 23075 6765 23076
rect 6270 23074 6336 23075
rect 6694 23074 6760 23075
rect 6270 22745 6336 22746
rect 6694 22745 6760 22746
rect 6265 22744 6271 22745
rect 5022 22733 5088 22734
rect 5494 22733 5560 22734
rect 5926 22733 5992 22734
rect 4980 22669 5023 22733
rect 5087 22669 5130 22733
rect 5452 22669 5495 22733
rect 5559 22669 5602 22733
rect 5884 22669 5927 22733
rect 5991 22669 6034 22733
rect 6228 22681 6271 22744
rect 6335 22744 6341 22745
rect 6689 22744 6695 22745
rect 6335 22681 6378 22744
rect 6228 22680 6378 22681
rect 6652 22681 6695 22744
rect 6759 22744 6765 22745
rect 6759 22681 6802 22744
rect 6652 22680 6802 22681
rect 5022 22668 5088 22669
rect 5494 22668 5560 22669
rect 5926 22668 5992 22669
rect 5022 22361 5088 22362
rect 5494 22361 5560 22362
rect 5926 22361 5992 22362
rect 4980 22297 5023 22361
rect 5087 22297 5130 22361
rect 5452 22297 5495 22361
rect 5559 22297 5602 22361
rect 5884 22297 5927 22361
rect 5991 22297 6034 22361
rect 6228 22349 6378 22350
rect 5022 22296 5088 22297
rect 5494 22296 5560 22297
rect 5926 22296 5992 22297
rect 6228 22286 6271 22349
rect 6265 22285 6271 22286
rect 6335 22286 6378 22349
rect 6652 22349 6802 22350
rect 6652 22286 6695 22349
rect 6335 22285 6341 22286
rect 6689 22285 6695 22286
rect 6759 22286 6802 22349
rect 6759 22285 6765 22286
rect 6270 22284 6336 22285
rect 6694 22284 6760 22285
rect 6270 21955 6336 21956
rect 6694 21955 6760 21956
rect 6265 21954 6271 21955
rect 5022 21943 5088 21944
rect 5494 21943 5560 21944
rect 5926 21943 5992 21944
rect 4980 21879 5023 21943
rect 5087 21879 5130 21943
rect 5452 21879 5495 21943
rect 5559 21879 5602 21943
rect 5884 21879 5927 21943
rect 5991 21879 6034 21943
rect 6228 21891 6271 21954
rect 6335 21954 6341 21955
rect 6689 21954 6695 21955
rect 6335 21891 6378 21954
rect 6228 21890 6378 21891
rect 6652 21891 6695 21954
rect 6759 21954 6765 21955
rect 6759 21891 6802 21954
rect 6652 21890 6802 21891
rect 5022 21878 5088 21879
rect 5494 21878 5560 21879
rect 5926 21878 5992 21879
rect 5022 21571 5088 21572
rect 5494 21571 5560 21572
rect 5926 21571 5992 21572
rect 4980 21507 5023 21571
rect 5087 21507 5130 21571
rect 5452 21507 5495 21571
rect 5559 21507 5602 21571
rect 5884 21507 5927 21571
rect 5991 21507 6034 21571
rect 6228 21559 6378 21560
rect 5022 21506 5088 21507
rect 5494 21506 5560 21507
rect 5926 21506 5992 21507
rect 6228 21496 6271 21559
rect 6265 21495 6271 21496
rect 6335 21496 6378 21559
rect 6652 21559 6802 21560
rect 6652 21496 6695 21559
rect 6335 21495 6341 21496
rect 6689 21495 6695 21496
rect 6759 21496 6802 21559
rect 6759 21495 6765 21496
rect 6270 21494 6336 21495
rect 6694 21494 6760 21495
rect 6270 21165 6336 21166
rect 6694 21165 6760 21166
rect 6265 21164 6271 21165
rect 5022 21153 5088 21154
rect 5494 21153 5560 21154
rect 5926 21153 5992 21154
rect 4980 21089 5023 21153
rect 5087 21089 5130 21153
rect 5452 21089 5495 21153
rect 5559 21089 5602 21153
rect 5884 21089 5927 21153
rect 5991 21089 6034 21153
rect 6228 21101 6271 21164
rect 6335 21164 6341 21165
rect 6689 21164 6695 21165
rect 6335 21101 6378 21164
rect 6228 21100 6378 21101
rect 6652 21101 6695 21164
rect 6759 21164 6765 21165
rect 6759 21101 6802 21164
rect 6652 21100 6802 21101
rect 5022 21088 5088 21089
rect 5494 21088 5560 21089
rect 5926 21088 5992 21089
rect 5022 20781 5088 20782
rect 5494 20781 5560 20782
rect 5926 20781 5992 20782
rect 4980 20717 5023 20781
rect 5087 20717 5130 20781
rect 5452 20717 5495 20781
rect 5559 20717 5602 20781
rect 5884 20717 5927 20781
rect 5991 20717 6034 20781
rect 6228 20769 6378 20770
rect 5022 20716 5088 20717
rect 5494 20716 5560 20717
rect 5926 20716 5992 20717
rect 6228 20706 6271 20769
rect 6265 20705 6271 20706
rect 6335 20706 6378 20769
rect 6652 20769 6802 20770
rect 6652 20706 6695 20769
rect 6335 20705 6341 20706
rect 6689 20705 6695 20706
rect 6759 20706 6802 20769
rect 6759 20705 6765 20706
rect 6270 20704 6336 20705
rect 6694 20704 6760 20705
rect 6270 20375 6336 20376
rect 6694 20375 6760 20376
rect 6265 20374 6271 20375
rect 5022 20363 5088 20364
rect 5494 20363 5560 20364
rect 5926 20363 5992 20364
rect 4980 20299 5023 20363
rect 5087 20299 5130 20363
rect 5452 20299 5495 20363
rect 5559 20299 5602 20363
rect 5884 20299 5927 20363
rect 5991 20299 6034 20363
rect 6228 20311 6271 20374
rect 6335 20374 6341 20375
rect 6689 20374 6695 20375
rect 6335 20311 6378 20374
rect 6228 20310 6378 20311
rect 6652 20311 6695 20374
rect 6759 20374 6765 20375
rect 6759 20311 6802 20374
rect 6652 20310 6802 20311
rect 5022 20298 5088 20299
rect 5494 20298 5560 20299
rect 5926 20298 5992 20299
rect 5022 19991 5088 19992
rect 5494 19991 5560 19992
rect 5926 19991 5992 19992
rect 4980 19927 5023 19991
rect 5087 19927 5130 19991
rect 5452 19927 5495 19991
rect 5559 19927 5602 19991
rect 5884 19927 5927 19991
rect 5991 19927 6034 19991
rect 6228 19979 6378 19980
rect 5022 19926 5088 19927
rect 5494 19926 5560 19927
rect 5926 19926 5992 19927
rect 6228 19916 6271 19979
rect 6265 19915 6271 19916
rect 6335 19916 6378 19979
rect 6652 19979 6802 19980
rect 6652 19916 6695 19979
rect 6335 19915 6341 19916
rect 6689 19915 6695 19916
rect 6759 19916 6802 19979
rect 6759 19915 6765 19916
rect 6270 19914 6336 19915
rect 6694 19914 6760 19915
rect 6270 19585 6336 19586
rect 6694 19585 6760 19586
rect 6265 19584 6271 19585
rect 5022 19573 5088 19574
rect 5494 19573 5560 19574
rect 5926 19573 5992 19574
rect 4980 19509 5023 19573
rect 5087 19509 5130 19573
rect 5452 19509 5495 19573
rect 5559 19509 5602 19573
rect 5884 19509 5927 19573
rect 5991 19509 6034 19573
rect 6228 19521 6271 19584
rect 6335 19584 6341 19585
rect 6689 19584 6695 19585
rect 6335 19521 6378 19584
rect 6228 19520 6378 19521
rect 6652 19521 6695 19584
rect 6759 19584 6765 19585
rect 6759 19521 6802 19584
rect 6652 19520 6802 19521
rect 5022 19508 5088 19509
rect 5494 19508 5560 19509
rect 5926 19508 5992 19509
rect 5022 19201 5088 19202
rect 5494 19201 5560 19202
rect 5926 19201 5992 19202
rect 4980 19137 5023 19201
rect 5087 19137 5130 19201
rect 5452 19137 5495 19201
rect 5559 19137 5602 19201
rect 5884 19137 5927 19201
rect 5991 19137 6034 19201
rect 6228 19189 6378 19190
rect 5022 19136 5088 19137
rect 5494 19136 5560 19137
rect 5926 19136 5992 19137
rect 6228 19126 6271 19189
rect 6265 19125 6271 19126
rect 6335 19126 6378 19189
rect 6652 19189 6802 19190
rect 6652 19126 6695 19189
rect 6335 19125 6341 19126
rect 6689 19125 6695 19126
rect 6759 19126 6802 19189
rect 6759 19125 6765 19126
rect 6270 19124 6336 19125
rect 6694 19124 6760 19125
rect 6270 18795 6336 18796
rect 6694 18795 6760 18796
rect 6265 18794 6271 18795
rect 5022 18783 5088 18784
rect 5494 18783 5560 18784
rect 5926 18783 5992 18784
rect 4980 18719 5023 18783
rect 5087 18719 5130 18783
rect 5452 18719 5495 18783
rect 5559 18719 5602 18783
rect 5884 18719 5927 18783
rect 5991 18719 6034 18783
rect 6228 18731 6271 18794
rect 6335 18794 6341 18795
rect 6689 18794 6695 18795
rect 6335 18731 6378 18794
rect 6228 18730 6378 18731
rect 6652 18731 6695 18794
rect 6759 18794 6765 18795
rect 6759 18731 6802 18794
rect 6652 18730 6802 18731
rect 5022 18718 5088 18719
rect 5494 18718 5560 18719
rect 5926 18718 5992 18719
rect 5022 18411 5088 18412
rect 5494 18411 5560 18412
rect 5926 18411 5992 18412
rect 4980 18347 5023 18411
rect 5087 18347 5130 18411
rect 5452 18347 5495 18411
rect 5559 18347 5602 18411
rect 5884 18347 5927 18411
rect 5991 18347 6034 18411
rect 6228 18399 6378 18400
rect 5022 18346 5088 18347
rect 5494 18346 5560 18347
rect 5926 18346 5992 18347
rect 6228 18336 6271 18399
rect 6265 18335 6271 18336
rect 6335 18336 6378 18399
rect 6652 18399 6802 18400
rect 6652 18336 6695 18399
rect 6335 18335 6341 18336
rect 6689 18335 6695 18336
rect 6759 18336 6802 18399
rect 6759 18335 6765 18336
rect 6270 18334 6336 18335
rect 6694 18334 6760 18335
rect 6270 18005 6336 18006
rect 6694 18005 6760 18006
rect 6265 18004 6271 18005
rect 5022 17993 5088 17994
rect 5494 17993 5560 17994
rect 5926 17993 5992 17994
rect 4980 17929 5023 17993
rect 5087 17929 5130 17993
rect 5452 17929 5495 17993
rect 5559 17929 5602 17993
rect 5884 17929 5927 17993
rect 5991 17929 6034 17993
rect 6228 17941 6271 18004
rect 6335 18004 6341 18005
rect 6689 18004 6695 18005
rect 6335 17941 6378 18004
rect 6228 17940 6378 17941
rect 6652 17941 6695 18004
rect 6759 18004 6765 18005
rect 6759 17941 6802 18004
rect 6652 17940 6802 17941
rect 5022 17928 5088 17929
rect 5494 17928 5560 17929
rect 5926 17928 5992 17929
rect 5022 17621 5088 17622
rect 5494 17621 5560 17622
rect 5926 17621 5992 17622
rect 4980 17557 5023 17621
rect 5087 17557 5130 17621
rect 5452 17557 5495 17621
rect 5559 17557 5602 17621
rect 5884 17557 5927 17621
rect 5991 17557 6034 17621
rect 6228 17609 6378 17610
rect 5022 17556 5088 17557
rect 5494 17556 5560 17557
rect 5926 17556 5992 17557
rect 6228 17546 6271 17609
rect 6265 17545 6271 17546
rect 6335 17546 6378 17609
rect 6652 17609 6802 17610
rect 6652 17546 6695 17609
rect 6335 17545 6341 17546
rect 6689 17545 6695 17546
rect 6759 17546 6802 17609
rect 6759 17545 6765 17546
rect 6270 17544 6336 17545
rect 6694 17544 6760 17545
rect 6270 17215 6336 17216
rect 6694 17215 6760 17216
rect 6265 17214 6271 17215
rect 5022 17203 5088 17204
rect 5494 17203 5560 17204
rect 5926 17203 5992 17204
rect 4980 17139 5023 17203
rect 5087 17139 5130 17203
rect 5452 17139 5495 17203
rect 5559 17139 5602 17203
rect 5884 17139 5927 17203
rect 5991 17139 6034 17203
rect 6228 17151 6271 17214
rect 6335 17214 6341 17215
rect 6689 17214 6695 17215
rect 6335 17151 6378 17214
rect 6228 17150 6378 17151
rect 6652 17151 6695 17214
rect 6759 17214 6765 17215
rect 6759 17151 6802 17214
rect 6652 17150 6802 17151
rect 5022 17138 5088 17139
rect 5494 17138 5560 17139
rect 5926 17138 5992 17139
rect 5022 16831 5088 16832
rect 5494 16831 5560 16832
rect 5926 16831 5992 16832
rect 4980 16767 5023 16831
rect 5087 16767 5130 16831
rect 5452 16767 5495 16831
rect 5559 16767 5602 16831
rect 5884 16767 5927 16831
rect 5991 16767 6034 16831
rect 6228 16819 6378 16820
rect 5022 16766 5088 16767
rect 5494 16766 5560 16767
rect 5926 16766 5992 16767
rect 6228 16756 6271 16819
rect 6265 16755 6271 16756
rect 6335 16756 6378 16819
rect 6652 16819 6802 16820
rect 6652 16756 6695 16819
rect 6335 16755 6341 16756
rect 6689 16755 6695 16756
rect 6759 16756 6802 16819
rect 6759 16755 6765 16756
rect 6270 16754 6336 16755
rect 6694 16754 6760 16755
rect 6270 16425 6336 16426
rect 6694 16425 6760 16426
rect 6265 16424 6271 16425
rect 5022 16413 5088 16414
rect 5494 16413 5560 16414
rect 5926 16413 5992 16414
rect 4980 16349 5023 16413
rect 5087 16349 5130 16413
rect 5452 16349 5495 16413
rect 5559 16349 5602 16413
rect 5884 16349 5927 16413
rect 5991 16349 6034 16413
rect 6228 16361 6271 16424
rect 6335 16424 6341 16425
rect 6689 16424 6695 16425
rect 6335 16361 6378 16424
rect 6228 16360 6378 16361
rect 6652 16361 6695 16424
rect 6759 16424 6765 16425
rect 6759 16361 6802 16424
rect 6652 16360 6802 16361
rect 5022 16348 5088 16349
rect 5494 16348 5560 16349
rect 5926 16348 5992 16349
rect 5022 16041 5088 16042
rect 5494 16041 5560 16042
rect 5926 16041 5992 16042
rect 4980 15977 5023 16041
rect 5087 15977 5130 16041
rect 5452 15977 5495 16041
rect 5559 15977 5602 16041
rect 5884 15977 5927 16041
rect 5991 15977 6034 16041
rect 6228 16029 6378 16030
rect 5022 15976 5088 15977
rect 5494 15976 5560 15977
rect 5926 15976 5992 15977
rect 6228 15966 6271 16029
rect 6265 15965 6271 15966
rect 6335 15966 6378 16029
rect 6652 16029 6802 16030
rect 6652 15966 6695 16029
rect 6335 15965 6341 15966
rect 6689 15965 6695 15966
rect 6759 15966 6802 16029
rect 6759 15965 6765 15966
rect 6270 15964 6336 15965
rect 6694 15964 6760 15965
rect 6270 15635 6336 15636
rect 6694 15635 6760 15636
rect 6265 15634 6271 15635
rect 5022 15623 5088 15624
rect 5494 15623 5560 15624
rect 5926 15623 5992 15624
rect 4980 15559 5023 15623
rect 5087 15559 5130 15623
rect 5452 15559 5495 15623
rect 5559 15559 5602 15623
rect 5884 15559 5927 15623
rect 5991 15559 6034 15623
rect 6228 15571 6271 15634
rect 6335 15634 6341 15635
rect 6689 15634 6695 15635
rect 6335 15571 6378 15634
rect 6228 15570 6378 15571
rect 6652 15571 6695 15634
rect 6759 15634 6765 15635
rect 6759 15571 6802 15634
rect 6652 15570 6802 15571
rect 5022 15558 5088 15559
rect 5494 15558 5560 15559
rect 5926 15558 5992 15559
rect 5022 15251 5088 15252
rect 5494 15251 5560 15252
rect 5926 15251 5992 15252
rect 4980 15187 5023 15251
rect 5087 15187 5130 15251
rect 5452 15187 5495 15251
rect 5559 15187 5602 15251
rect 5884 15187 5927 15251
rect 5991 15187 6034 15251
rect 6228 15239 6378 15240
rect 5022 15186 5088 15187
rect 5494 15186 5560 15187
rect 5926 15186 5992 15187
rect 6228 15176 6271 15239
rect 6265 15175 6271 15176
rect 6335 15176 6378 15239
rect 6652 15239 6802 15240
rect 6652 15176 6695 15239
rect 6335 15175 6341 15176
rect 6689 15175 6695 15176
rect 6759 15176 6802 15239
rect 6759 15175 6765 15176
rect 6270 15174 6336 15175
rect 6694 15174 6760 15175
rect 6270 14845 6336 14846
rect 6694 14845 6760 14846
rect 6265 14844 6271 14845
rect 5022 14833 5088 14834
rect 5494 14833 5560 14834
rect 5926 14833 5992 14834
rect 4980 14769 5023 14833
rect 5087 14769 5130 14833
rect 5452 14769 5495 14833
rect 5559 14769 5602 14833
rect 5884 14769 5927 14833
rect 5991 14769 6034 14833
rect 6228 14781 6271 14844
rect 6335 14844 6341 14845
rect 6689 14844 6695 14845
rect 6335 14781 6378 14844
rect 6228 14780 6378 14781
rect 6652 14781 6695 14844
rect 6759 14844 6765 14845
rect 6759 14781 6802 14844
rect 6652 14780 6802 14781
rect 5022 14768 5088 14769
rect 5494 14768 5560 14769
rect 5926 14768 5992 14769
rect 5022 14461 5088 14462
rect 5494 14461 5560 14462
rect 5926 14461 5992 14462
rect 4980 14397 5023 14461
rect 5087 14397 5130 14461
rect 5452 14397 5495 14461
rect 5559 14397 5602 14461
rect 5884 14397 5927 14461
rect 5991 14397 6034 14461
rect 6228 14449 6378 14450
rect 5022 14396 5088 14397
rect 5494 14396 5560 14397
rect 5926 14396 5992 14397
rect 6228 14386 6271 14449
rect 6265 14385 6271 14386
rect 6335 14386 6378 14449
rect 6652 14449 6802 14450
rect 6652 14386 6695 14449
rect 6335 14385 6341 14386
rect 6689 14385 6695 14386
rect 6759 14386 6802 14449
rect 6759 14385 6765 14386
rect 6270 14384 6336 14385
rect 6694 14384 6760 14385
rect 6270 14055 6336 14056
rect 6694 14055 6760 14056
rect 6265 14054 6271 14055
rect 5022 14043 5088 14044
rect 5494 14043 5560 14044
rect 5926 14043 5992 14044
rect 4980 13979 5023 14043
rect 5087 13979 5130 14043
rect 5452 13979 5495 14043
rect 5559 13979 5602 14043
rect 5884 13979 5927 14043
rect 5991 13979 6034 14043
rect 6228 13991 6271 14054
rect 6335 14054 6341 14055
rect 6689 14054 6695 14055
rect 6335 13991 6378 14054
rect 6228 13990 6378 13991
rect 6652 13991 6695 14054
rect 6759 14054 6765 14055
rect 6759 13991 6802 14054
rect 6652 13990 6802 13991
rect 5022 13978 5088 13979
rect 5494 13978 5560 13979
rect 5926 13978 5992 13979
rect 5022 13671 5088 13672
rect 5494 13671 5560 13672
rect 5926 13671 5992 13672
rect 4980 13607 5023 13671
rect 5087 13607 5130 13671
rect 5452 13607 5495 13671
rect 5559 13607 5602 13671
rect 5884 13607 5927 13671
rect 5991 13607 6034 13671
rect 6228 13659 6378 13660
rect 5022 13606 5088 13607
rect 5494 13606 5560 13607
rect 5926 13606 5992 13607
rect 6228 13596 6271 13659
rect 6265 13595 6271 13596
rect 6335 13596 6378 13659
rect 6652 13659 6802 13660
rect 6652 13596 6695 13659
rect 6335 13595 6341 13596
rect 6689 13595 6695 13596
rect 6759 13596 6802 13659
rect 6759 13595 6765 13596
rect 6270 13594 6336 13595
rect 6694 13594 6760 13595
rect 6270 13265 6336 13266
rect 6694 13265 6760 13266
rect 6265 13264 6271 13265
rect 5022 13253 5088 13254
rect 5494 13253 5560 13254
rect 5926 13253 5992 13254
rect 4980 13189 5023 13253
rect 5087 13189 5130 13253
rect 5452 13189 5495 13253
rect 5559 13189 5602 13253
rect 5884 13189 5927 13253
rect 5991 13189 6034 13253
rect 6228 13201 6271 13264
rect 6335 13264 6341 13265
rect 6689 13264 6695 13265
rect 6335 13201 6378 13264
rect 6228 13200 6378 13201
rect 6652 13201 6695 13264
rect 6759 13264 6765 13265
rect 6759 13201 6802 13264
rect 6652 13200 6802 13201
rect 5022 13188 5088 13189
rect 5494 13188 5560 13189
rect 5926 13188 5992 13189
rect 5022 12881 5088 12882
rect 5494 12881 5560 12882
rect 5926 12881 5992 12882
rect 4980 12817 5023 12881
rect 5087 12817 5130 12881
rect 5452 12817 5495 12881
rect 5559 12817 5602 12881
rect 5884 12817 5927 12881
rect 5991 12817 6034 12881
rect 6228 12869 6378 12870
rect 5022 12816 5088 12817
rect 5494 12816 5560 12817
rect 5926 12816 5992 12817
rect 6228 12806 6271 12869
rect 6265 12805 6271 12806
rect 6335 12806 6378 12869
rect 6652 12869 6802 12870
rect 6652 12806 6695 12869
rect 6335 12805 6341 12806
rect 6689 12805 6695 12806
rect 6759 12806 6802 12869
rect 6759 12805 6765 12806
rect 6270 12804 6336 12805
rect 6694 12804 6760 12805
rect 6270 12475 6336 12476
rect 6694 12475 6760 12476
rect 6265 12474 6271 12475
rect 5022 12463 5088 12464
rect 5494 12463 5560 12464
rect 5926 12463 5992 12464
rect 4980 12399 5023 12463
rect 5087 12399 5130 12463
rect 5452 12399 5495 12463
rect 5559 12399 5602 12463
rect 5884 12399 5927 12463
rect 5991 12399 6034 12463
rect 6228 12411 6271 12474
rect 6335 12474 6341 12475
rect 6689 12474 6695 12475
rect 6335 12411 6378 12474
rect 6228 12410 6378 12411
rect 6652 12411 6695 12474
rect 6759 12474 6765 12475
rect 6759 12411 6802 12474
rect 6652 12410 6802 12411
rect 5022 12398 5088 12399
rect 5494 12398 5560 12399
rect 5926 12398 5992 12399
rect 5022 12091 5088 12092
rect 5494 12091 5560 12092
rect 5926 12091 5992 12092
rect 4980 12027 5023 12091
rect 5087 12027 5130 12091
rect 5452 12027 5495 12091
rect 5559 12027 5602 12091
rect 5884 12027 5927 12091
rect 5991 12027 6034 12091
rect 6228 12079 6378 12080
rect 5022 12026 5088 12027
rect 5494 12026 5560 12027
rect 5926 12026 5992 12027
rect 6228 12016 6271 12079
rect 6265 12015 6271 12016
rect 6335 12016 6378 12079
rect 6652 12079 6802 12080
rect 6652 12016 6695 12079
rect 6335 12015 6341 12016
rect 6689 12015 6695 12016
rect 6759 12016 6802 12079
rect 6759 12015 6765 12016
rect 6270 12014 6336 12015
rect 6694 12014 6760 12015
rect 6270 11685 6336 11686
rect 6694 11685 6760 11686
rect 6265 11684 6271 11685
rect 5022 11673 5088 11674
rect 5494 11673 5560 11674
rect 5926 11673 5992 11674
rect 4980 11609 5023 11673
rect 5087 11609 5130 11673
rect 5452 11609 5495 11673
rect 5559 11609 5602 11673
rect 5884 11609 5927 11673
rect 5991 11609 6034 11673
rect 6228 11621 6271 11684
rect 6335 11684 6341 11685
rect 6689 11684 6695 11685
rect 6335 11621 6378 11684
rect 6228 11620 6378 11621
rect 6652 11621 6695 11684
rect 6759 11684 6765 11685
rect 6759 11621 6802 11684
rect 6652 11620 6802 11621
rect 5022 11608 5088 11609
rect 5494 11608 5560 11609
rect 5926 11608 5992 11609
rect 5022 11301 5088 11302
rect 5494 11301 5560 11302
rect 5926 11301 5992 11302
rect 4980 11237 5023 11301
rect 5087 11237 5130 11301
rect 5452 11237 5495 11301
rect 5559 11237 5602 11301
rect 5884 11237 5927 11301
rect 5991 11237 6034 11301
rect 6228 11289 6378 11290
rect 5022 11236 5088 11237
rect 5494 11236 5560 11237
rect 5926 11236 5992 11237
rect 6228 11226 6271 11289
rect 6265 11225 6271 11226
rect 6335 11226 6378 11289
rect 6652 11289 6802 11290
rect 6652 11226 6695 11289
rect 6335 11225 6341 11226
rect 6689 11225 6695 11226
rect 6759 11226 6802 11289
rect 6759 11225 6765 11226
rect 6270 11224 6336 11225
rect 6694 11224 6760 11225
rect 6270 10895 6336 10896
rect 6694 10895 6760 10896
rect 6265 10894 6271 10895
rect 5022 10883 5088 10884
rect 5494 10883 5560 10884
rect 5926 10883 5992 10884
rect 4980 10819 5023 10883
rect 5087 10819 5130 10883
rect 5452 10819 5495 10883
rect 5559 10819 5602 10883
rect 5884 10819 5927 10883
rect 5991 10819 6034 10883
rect 6228 10831 6271 10894
rect 6335 10894 6341 10895
rect 6689 10894 6695 10895
rect 6335 10831 6378 10894
rect 6228 10830 6378 10831
rect 6652 10831 6695 10894
rect 6759 10894 6765 10895
rect 6759 10831 6802 10894
rect 6652 10830 6802 10831
rect 5022 10818 5088 10819
rect 5494 10818 5560 10819
rect 5926 10818 5992 10819
rect 5022 10511 5088 10512
rect 5494 10511 5560 10512
rect 5926 10511 5992 10512
rect 4980 10447 5023 10511
rect 5087 10447 5130 10511
rect 5452 10447 5495 10511
rect 5559 10447 5602 10511
rect 5884 10447 5927 10511
rect 5991 10447 6034 10511
rect 6228 10499 6378 10500
rect 5022 10446 5088 10447
rect 5494 10446 5560 10447
rect 5926 10446 5992 10447
rect 6228 10436 6271 10499
rect 6265 10435 6271 10436
rect 6335 10436 6378 10499
rect 6652 10499 6802 10500
rect 6652 10436 6695 10499
rect 6335 10435 6341 10436
rect 6689 10435 6695 10436
rect 6759 10436 6802 10499
rect 6759 10435 6765 10436
rect 6270 10434 6336 10435
rect 6694 10434 6760 10435
rect 6270 10105 6336 10106
rect 6694 10105 6760 10106
rect 6265 10104 6271 10105
rect 5022 10093 5088 10094
rect 5494 10093 5560 10094
rect 5926 10093 5992 10094
rect 4980 10029 5023 10093
rect 5087 10029 5130 10093
rect 5452 10029 5495 10093
rect 5559 10029 5602 10093
rect 5884 10029 5927 10093
rect 5991 10029 6034 10093
rect 6228 10041 6271 10104
rect 6335 10104 6341 10105
rect 6689 10104 6695 10105
rect 6335 10041 6378 10104
rect 6228 10040 6378 10041
rect 6652 10041 6695 10104
rect 6759 10104 6765 10105
rect 6759 10041 6802 10104
rect 6652 10040 6802 10041
rect 5022 10028 5088 10029
rect 5494 10028 5560 10029
rect 5926 10028 5992 10029
rect 5022 9721 5088 9722
rect 5494 9721 5560 9722
rect 5926 9721 5992 9722
rect 4980 9657 5023 9721
rect 5087 9657 5130 9721
rect 5452 9657 5495 9721
rect 5559 9657 5602 9721
rect 5884 9657 5927 9721
rect 5991 9657 6034 9721
rect 6228 9709 6378 9710
rect 5022 9656 5088 9657
rect 5494 9656 5560 9657
rect 5926 9656 5992 9657
rect 6228 9646 6271 9709
rect 6265 9645 6271 9646
rect 6335 9646 6378 9709
rect 6652 9709 6802 9710
rect 6652 9646 6695 9709
rect 6335 9645 6341 9646
rect 6689 9645 6695 9646
rect 6759 9646 6802 9709
rect 6759 9645 6765 9646
rect 6270 9644 6336 9645
rect 6694 9644 6760 9645
rect 6270 9315 6336 9316
rect 6694 9315 6760 9316
rect 6265 9314 6271 9315
rect 5022 9303 5088 9304
rect 5494 9303 5560 9304
rect 5926 9303 5992 9304
rect 4980 9239 5023 9303
rect 5087 9239 5130 9303
rect 5452 9239 5495 9303
rect 5559 9239 5602 9303
rect 5884 9239 5927 9303
rect 5991 9239 6034 9303
rect 6228 9251 6271 9314
rect 6335 9314 6341 9315
rect 6689 9314 6695 9315
rect 6335 9251 6378 9314
rect 6228 9250 6378 9251
rect 6652 9251 6695 9314
rect 6759 9314 6765 9315
rect 6759 9251 6802 9314
rect 6652 9250 6802 9251
rect 5022 9238 5088 9239
rect 5494 9238 5560 9239
rect 5926 9238 5992 9239
rect 5022 8931 5088 8932
rect 5494 8931 5560 8932
rect 5926 8931 5992 8932
rect 4980 8867 5023 8931
rect 5087 8867 5130 8931
rect 5452 8867 5495 8931
rect 5559 8867 5602 8931
rect 5884 8867 5927 8931
rect 5991 8867 6034 8931
rect 6228 8919 6378 8920
rect 5022 8866 5088 8867
rect 5494 8866 5560 8867
rect 5926 8866 5992 8867
rect 6228 8856 6271 8919
rect 6265 8855 6271 8856
rect 6335 8856 6378 8919
rect 6652 8919 6802 8920
rect 6652 8856 6695 8919
rect 6335 8855 6341 8856
rect 6689 8855 6695 8856
rect 6759 8856 6802 8919
rect 6759 8855 6765 8856
rect 6270 8854 6336 8855
rect 6694 8854 6760 8855
rect 6270 8525 6336 8526
rect 6694 8525 6760 8526
rect 6265 8524 6271 8525
rect 5022 8513 5088 8514
rect 5494 8513 5560 8514
rect 5926 8513 5992 8514
rect 4980 8449 5023 8513
rect 5087 8449 5130 8513
rect 5452 8449 5495 8513
rect 5559 8449 5602 8513
rect 5884 8449 5927 8513
rect 5991 8449 6034 8513
rect 6228 8461 6271 8524
rect 6335 8524 6341 8525
rect 6689 8524 6695 8525
rect 6335 8461 6378 8524
rect 6228 8460 6378 8461
rect 6652 8461 6695 8524
rect 6759 8524 6765 8525
rect 6759 8461 6802 8524
rect 6652 8460 6802 8461
rect 5022 8448 5088 8449
rect 5494 8448 5560 8449
rect 5926 8448 5992 8449
rect 5022 8141 5088 8142
rect 5494 8141 5560 8142
rect 5926 8141 5992 8142
rect 4980 8077 5023 8141
rect 5087 8077 5130 8141
rect 5452 8077 5495 8141
rect 5559 8077 5602 8141
rect 5884 8077 5927 8141
rect 5991 8077 6034 8141
rect 6228 8129 6378 8130
rect 5022 8076 5088 8077
rect 5494 8076 5560 8077
rect 5926 8076 5992 8077
rect 6228 8066 6271 8129
rect 6265 8065 6271 8066
rect 6335 8066 6378 8129
rect 6652 8129 6802 8130
rect 6652 8066 6695 8129
rect 6335 8065 6341 8066
rect 6689 8065 6695 8066
rect 6759 8066 6802 8129
rect 6759 8065 6765 8066
rect 6270 8064 6336 8065
rect 6694 8064 6760 8065
rect 6270 7735 6336 7736
rect 6694 7735 6760 7736
rect 6265 7734 6271 7735
rect 5022 7723 5088 7724
rect 5494 7723 5560 7724
rect 5926 7723 5992 7724
rect 4980 7659 5023 7723
rect 5087 7659 5130 7723
rect 5452 7659 5495 7723
rect 5559 7659 5602 7723
rect 5884 7659 5927 7723
rect 5991 7659 6034 7723
rect 6228 7671 6271 7734
rect 6335 7734 6341 7735
rect 6689 7734 6695 7735
rect 6335 7671 6378 7734
rect 6228 7670 6378 7671
rect 6652 7671 6695 7734
rect 6759 7734 6765 7735
rect 6759 7671 6802 7734
rect 6652 7670 6802 7671
rect 5022 7658 5088 7659
rect 5494 7658 5560 7659
rect 5926 7658 5992 7659
rect 5022 7351 5088 7352
rect 5494 7351 5560 7352
rect 5926 7351 5992 7352
rect 4980 7287 5023 7351
rect 5087 7287 5130 7351
rect 5452 7287 5495 7351
rect 5559 7287 5602 7351
rect 5884 7287 5927 7351
rect 5991 7287 6034 7351
rect 6228 7339 6378 7340
rect 5022 7286 5088 7287
rect 5494 7286 5560 7287
rect 5926 7286 5992 7287
rect 6228 7276 6271 7339
rect 6265 7275 6271 7276
rect 6335 7276 6378 7339
rect 6652 7339 6802 7340
rect 6652 7276 6695 7339
rect 6335 7275 6341 7276
rect 6689 7275 6695 7276
rect 6759 7276 6802 7339
rect 6759 7275 6765 7276
rect 6270 7274 6336 7275
rect 6694 7274 6760 7275
rect 6270 6945 6336 6946
rect 6694 6945 6760 6946
rect 6265 6944 6271 6945
rect 5022 6933 5088 6934
rect 5494 6933 5560 6934
rect 5926 6933 5992 6934
rect 4980 6869 5023 6933
rect 5087 6869 5130 6933
rect 5452 6869 5495 6933
rect 5559 6869 5602 6933
rect 5884 6869 5927 6933
rect 5991 6869 6034 6933
rect 6228 6881 6271 6944
rect 6335 6944 6341 6945
rect 6689 6944 6695 6945
rect 6335 6881 6378 6944
rect 6228 6880 6378 6881
rect 6652 6881 6695 6944
rect 6759 6944 6765 6945
rect 6759 6881 6802 6944
rect 6652 6880 6802 6881
rect 5022 6868 5088 6869
rect 5494 6868 5560 6869
rect 5926 6868 5992 6869
rect 5022 6561 5088 6562
rect 5494 6561 5560 6562
rect 5926 6561 5992 6562
rect 4980 6497 5023 6561
rect 5087 6497 5130 6561
rect 5452 6497 5495 6561
rect 5559 6497 5602 6561
rect 5884 6497 5927 6561
rect 5991 6497 6034 6561
rect 6228 6549 6378 6550
rect 5022 6496 5088 6497
rect 5494 6496 5560 6497
rect 5926 6496 5992 6497
rect 6228 6486 6271 6549
rect 6265 6485 6271 6486
rect 6335 6486 6378 6549
rect 6652 6549 6802 6550
rect 6652 6486 6695 6549
rect 6335 6485 6341 6486
rect 6689 6485 6695 6486
rect 6759 6486 6802 6549
rect 6759 6485 6765 6486
rect 6270 6484 6336 6485
rect 6694 6484 6760 6485
rect 6270 6155 6336 6156
rect 6694 6155 6760 6156
rect 6265 6154 6271 6155
rect 5022 6143 5088 6144
rect 5494 6143 5560 6144
rect 5926 6143 5992 6144
rect 4980 6079 5023 6143
rect 5087 6079 5130 6143
rect 5452 6079 5495 6143
rect 5559 6079 5602 6143
rect 5884 6079 5927 6143
rect 5991 6079 6034 6143
rect 6228 6091 6271 6154
rect 6335 6154 6341 6155
rect 6689 6154 6695 6155
rect 6335 6091 6378 6154
rect 6228 6090 6378 6091
rect 6652 6091 6695 6154
rect 6759 6154 6765 6155
rect 6759 6091 6802 6154
rect 6652 6090 6802 6091
rect 5022 6078 5088 6079
rect 5494 6078 5560 6079
rect 5926 6078 5992 6079
rect 2290 5883 2388 5981
rect 2715 5883 2813 5981
rect 3094 5876 3192 5974
rect 3490 5876 3588 5974
rect 5022 5771 5088 5772
rect 5494 5771 5560 5772
rect 5926 5771 5992 5772
rect 4980 5707 5023 5771
rect 5087 5707 5130 5771
rect 5452 5707 5495 5771
rect 5559 5707 5602 5771
rect 5884 5707 5927 5771
rect 5991 5707 6034 5771
rect 6228 5759 6378 5760
rect 5022 5706 5088 5707
rect 5494 5706 5560 5707
rect 5926 5706 5992 5707
rect 6228 5696 6271 5759
rect 6265 5695 6271 5696
rect 6335 5696 6378 5759
rect 6652 5759 6802 5760
rect 6652 5696 6695 5759
rect 6335 5695 6341 5696
rect 6689 5695 6695 5696
rect 6759 5696 6802 5759
rect 6759 5695 6765 5696
rect 6270 5694 6336 5695
rect 6694 5694 6760 5695
rect 6270 5365 6336 5366
rect 6694 5365 6760 5366
rect 6265 5364 6271 5365
rect 5022 5353 5088 5354
rect 5494 5353 5560 5354
rect 5926 5353 5992 5354
rect 4980 5289 5023 5353
rect 5087 5289 5130 5353
rect 5452 5289 5495 5353
rect 5559 5289 5602 5353
rect 5884 5289 5927 5353
rect 5991 5289 6034 5353
rect 6228 5301 6271 5364
rect 6335 5364 6341 5365
rect 6689 5364 6695 5365
rect 6335 5301 6378 5364
rect 6228 5300 6378 5301
rect 6652 5301 6695 5364
rect 6759 5364 6765 5365
rect 6759 5301 6802 5364
rect 6652 5300 6802 5301
rect 5022 5288 5088 5289
rect 5494 5288 5560 5289
rect 5926 5288 5992 5289
rect 996 5086 1094 5184
rect 1392 5086 1490 5184
rect 2290 5093 2388 5191
rect 2715 5093 2813 5191
rect 3094 5086 3192 5184
rect 3490 5086 3588 5184
rect 5022 4981 5088 4982
rect 5494 4981 5560 4982
rect 5926 4981 5992 4982
rect 4980 4917 5023 4981
rect 5087 4917 5130 4981
rect 5452 4917 5495 4981
rect 5559 4917 5602 4981
rect 5884 4917 5927 4981
rect 5991 4917 6034 4981
rect 6228 4969 6378 4970
rect 5022 4916 5088 4917
rect 5494 4916 5560 4917
rect 5926 4916 5992 4917
rect 6228 4906 6271 4969
rect 6265 4905 6271 4906
rect 6335 4906 6378 4969
rect 6652 4969 6802 4970
rect 6652 4906 6695 4969
rect 6335 4905 6341 4906
rect 6689 4905 6695 4906
rect 6759 4906 6802 4969
rect 6759 4905 6765 4906
rect 6270 4904 6336 4905
rect 6694 4904 6760 4905
rect 6270 4575 6336 4576
rect 6694 4575 6760 4576
rect 6265 4574 6271 4575
rect 5022 4563 5088 4564
rect 5494 4563 5560 4564
rect 5926 4563 5992 4564
rect 4980 4499 5023 4563
rect 5087 4499 5130 4563
rect 5452 4499 5495 4563
rect 5559 4499 5602 4563
rect 5884 4499 5927 4563
rect 5991 4499 6034 4563
rect 6228 4511 6271 4574
rect 6335 4574 6341 4575
rect 6689 4574 6695 4575
rect 6335 4511 6378 4574
rect 6228 4510 6378 4511
rect 6652 4511 6695 4574
rect 6759 4574 6765 4575
rect 6759 4511 6802 4574
rect 6652 4510 6802 4511
rect 5022 4498 5088 4499
rect 5494 4498 5560 4499
rect 5926 4498 5992 4499
rect 5022 4191 5088 4192
rect 5494 4191 5560 4192
rect 5926 4191 5992 4192
rect 4980 4127 5023 4191
rect 5087 4127 5130 4191
rect 5452 4127 5495 4191
rect 5559 4127 5602 4191
rect 5884 4127 5927 4191
rect 5991 4127 6034 4191
rect 6228 4179 6378 4180
rect 5022 4126 5088 4127
rect 5494 4126 5560 4127
rect 5926 4126 5992 4127
rect 6228 4116 6271 4179
rect 6265 4115 6271 4116
rect 6335 4116 6378 4179
rect 6652 4179 6802 4180
rect 6652 4116 6695 4179
rect 6335 4115 6341 4116
rect 6689 4115 6695 4116
rect 6759 4116 6802 4179
rect 6759 4115 6765 4116
rect 6270 4114 6336 4115
rect 6694 4114 6760 4115
rect 6270 3785 6336 3786
rect 6694 3785 6760 3786
rect 6265 3784 6271 3785
rect 5022 3773 5088 3774
rect 5494 3773 5560 3774
rect 5926 3773 5992 3774
rect 4980 3709 5023 3773
rect 5087 3709 5130 3773
rect 5452 3709 5495 3773
rect 5559 3709 5602 3773
rect 5884 3709 5927 3773
rect 5991 3709 6034 3773
rect 6228 3721 6271 3784
rect 6335 3784 6341 3785
rect 6689 3784 6695 3785
rect 6335 3721 6378 3784
rect 6228 3720 6378 3721
rect 6652 3721 6695 3784
rect 6759 3784 6765 3785
rect 6759 3721 6802 3784
rect 6652 3720 6802 3721
rect 5022 3708 5088 3709
rect 5494 3708 5560 3709
rect 5926 3708 5992 3709
rect 2290 3513 2388 3611
rect 2715 3513 2813 3611
rect 3094 3506 3192 3604
rect 3490 3506 3588 3604
rect 5022 3401 5088 3402
rect 5494 3401 5560 3402
rect 5926 3401 5992 3402
rect 4980 3337 5023 3401
rect 5087 3337 5130 3401
rect 5452 3337 5495 3401
rect 5559 3337 5602 3401
rect 5884 3337 5927 3401
rect 5991 3337 6034 3401
rect 6228 3389 6378 3390
rect 5022 3336 5088 3337
rect 5494 3336 5560 3337
rect 5926 3336 5992 3337
rect 6228 3326 6271 3389
rect 6265 3325 6271 3326
rect 6335 3326 6378 3389
rect 6652 3389 6802 3390
rect 6652 3326 6695 3389
rect 6335 3325 6341 3326
rect 6689 3325 6695 3326
rect 6759 3326 6802 3389
rect 6759 3325 6765 3326
rect 6270 3324 6336 3325
rect 6694 3324 6760 3325
rect 6270 2995 6336 2996
rect 6694 2995 6760 2996
rect 6265 2994 6271 2995
rect 5022 2983 5088 2984
rect 5494 2983 5560 2984
rect 5926 2983 5992 2984
rect 4980 2919 5023 2983
rect 5087 2919 5130 2983
rect 5452 2919 5495 2983
rect 5559 2919 5602 2983
rect 5884 2919 5927 2983
rect 5991 2919 6034 2983
rect 6228 2931 6271 2994
rect 6335 2994 6341 2995
rect 6689 2994 6695 2995
rect 6335 2931 6378 2994
rect 6228 2930 6378 2931
rect 6652 2931 6695 2994
rect 6759 2994 6765 2995
rect 6759 2931 6802 2994
rect 6652 2930 6802 2931
rect 5022 2918 5088 2919
rect 5494 2918 5560 2919
rect 5926 2918 5992 2919
rect 996 2716 1094 2814
rect 1392 2716 1490 2814
rect 2290 2723 2388 2821
rect 2715 2723 2813 2821
rect 3094 2716 3192 2814
rect 3490 2716 3588 2814
rect 5022 2611 5088 2612
rect 5494 2611 5560 2612
rect 5926 2611 5992 2612
rect 4980 2547 5023 2611
rect 5087 2547 5130 2611
rect 5452 2547 5495 2611
rect 5559 2547 5602 2611
rect 5884 2547 5927 2611
rect 5991 2547 6034 2611
rect 6228 2599 6378 2600
rect 5022 2546 5088 2547
rect 5494 2546 5560 2547
rect 5926 2546 5992 2547
rect 6228 2536 6271 2599
rect 6265 2535 6271 2536
rect 6335 2536 6378 2599
rect 6652 2599 6802 2600
rect 6652 2536 6695 2599
rect 6335 2535 6341 2536
rect 6689 2535 6695 2536
rect 6759 2536 6802 2599
rect 6759 2535 6765 2536
rect 6270 2534 6336 2535
rect 6694 2534 6760 2535
rect 6270 2205 6336 2206
rect 6694 2205 6760 2206
rect 6265 2204 6271 2205
rect 5022 2193 5088 2194
rect 5494 2193 5560 2194
rect 5926 2193 5992 2194
rect 4980 2129 5023 2193
rect 5087 2129 5130 2193
rect 5452 2129 5495 2193
rect 5559 2129 5602 2193
rect 5884 2129 5927 2193
rect 5991 2129 6034 2193
rect 6228 2141 6271 2204
rect 6335 2204 6341 2205
rect 6689 2204 6695 2205
rect 6335 2141 6378 2204
rect 6228 2140 6378 2141
rect 6652 2141 6695 2204
rect 6759 2204 6765 2205
rect 6759 2141 6802 2204
rect 6652 2140 6802 2141
rect 5022 2128 5088 2129
rect 5494 2128 5560 2129
rect 5926 2128 5992 2129
rect 5022 1821 5088 1822
rect 5494 1821 5560 1822
rect 5926 1821 5992 1822
rect 4980 1757 5023 1821
rect 5087 1757 5130 1821
rect 5452 1757 5495 1821
rect 5559 1757 5602 1821
rect 5884 1757 5927 1821
rect 5991 1757 6034 1821
rect 6228 1809 6378 1810
rect 5022 1756 5088 1757
rect 5494 1756 5560 1757
rect 5926 1756 5992 1757
rect 6228 1746 6271 1809
rect 6265 1745 6271 1746
rect 6335 1746 6378 1809
rect 6652 1809 6802 1810
rect 6652 1746 6695 1809
rect 6335 1745 6341 1746
rect 6689 1745 6695 1746
rect 6759 1746 6802 1809
rect 6759 1745 6765 1746
rect 6270 1744 6336 1745
rect 6694 1744 6760 1745
rect 6270 1415 6336 1416
rect 6694 1415 6760 1416
rect 6265 1414 6271 1415
rect 5022 1403 5088 1404
rect 5494 1403 5560 1404
rect 5926 1403 5992 1404
rect 4980 1339 5023 1403
rect 5087 1339 5130 1403
rect 5452 1339 5495 1403
rect 5559 1339 5602 1403
rect 5884 1339 5927 1403
rect 5991 1339 6034 1403
rect 6228 1351 6271 1414
rect 6335 1414 6341 1415
rect 6689 1414 6695 1415
rect 6335 1351 6378 1414
rect 6228 1350 6378 1351
rect 6652 1351 6695 1414
rect 6759 1414 6765 1415
rect 6759 1351 6802 1414
rect 6652 1350 6802 1351
rect 5022 1338 5088 1339
rect 5494 1338 5560 1339
rect 5926 1338 5992 1339
rect 2290 1143 2388 1241
rect 2715 1143 2813 1241
rect 3094 1136 3192 1234
rect 3490 1136 3588 1234
rect 5022 1031 5088 1032
rect 5494 1031 5560 1032
rect 5926 1031 5992 1032
rect 4980 967 5023 1031
rect 5087 967 5130 1031
rect 5452 967 5495 1031
rect 5559 967 5602 1031
rect 5884 967 5927 1031
rect 5991 967 6034 1031
rect 6228 1019 6378 1020
rect 5022 966 5088 967
rect 5494 966 5560 967
rect 5926 966 5992 967
rect 6228 956 6271 1019
rect 6265 955 6271 956
rect 6335 956 6378 1019
rect 6652 1019 6802 1020
rect 6652 956 6695 1019
rect 6335 955 6341 956
rect 6689 955 6695 956
rect 6759 956 6802 1019
rect 6759 955 6765 956
rect 6270 954 6336 955
rect 6694 954 6760 955
rect 6270 625 6336 626
rect 6694 625 6760 626
rect 6265 624 6271 625
rect 5022 613 5088 614
rect 5494 613 5560 614
rect 5926 613 5992 614
rect 4980 549 5023 613
rect 5087 549 5130 613
rect 5452 549 5495 613
rect 5559 549 5602 613
rect 5884 549 5927 613
rect 5991 549 6034 613
rect 6228 561 6271 624
rect 6335 624 6341 625
rect 6689 624 6695 625
rect 6335 561 6378 624
rect 6228 560 6378 561
rect 6652 561 6695 624
rect 6759 624 6765 625
rect 6759 561 6802 624
rect 6652 560 6802 561
rect 5022 548 5088 549
rect 5494 548 5560 549
rect 5926 548 5992 549
rect 996 346 1094 444
rect 1392 346 1490 444
rect 2290 353 2388 451
rect 2715 353 2813 451
rect 3094 346 3192 444
rect 3490 346 3588 444
rect 5022 241 5088 242
rect 5494 241 5560 242
rect 5926 241 5992 242
rect 4980 177 5023 241
rect 5087 177 5130 241
rect 5452 177 5495 241
rect 5559 177 5602 241
rect 5884 177 5927 241
rect 5991 177 6034 241
rect 6228 229 6378 230
rect 5022 176 5088 177
rect 5494 176 5560 177
rect 5926 176 5992 177
rect 6228 166 6271 229
rect 6265 165 6271 166
rect 6335 166 6378 229
rect 6652 229 6802 230
rect 6652 166 6695 229
rect 6335 165 6341 166
rect 6689 165 6695 166
rect 6759 166 6802 229
rect 6759 165 6765 166
rect 6270 164 6336 165
rect 6694 164 6760 165
<< via3 >>
rect 5023 25099 5087 25103
rect 5023 25043 5027 25099
rect 5027 25043 5083 25099
rect 5083 25043 5087 25099
rect 5023 25039 5087 25043
rect 5495 25099 5559 25103
rect 5495 25043 5499 25099
rect 5499 25043 5555 25099
rect 5555 25043 5559 25099
rect 5495 25039 5559 25043
rect 5927 25099 5991 25103
rect 5927 25043 5931 25099
rect 5931 25043 5987 25099
rect 5987 25043 5991 25099
rect 5927 25039 5991 25043
rect 6271 25111 6335 25115
rect 6271 25055 6275 25111
rect 6275 25055 6331 25111
rect 6331 25055 6335 25111
rect 6271 25051 6335 25055
rect 6695 25111 6759 25115
rect 6695 25055 6699 25111
rect 6699 25055 6755 25111
rect 6755 25055 6759 25111
rect 6695 25051 6759 25055
rect 5023 24727 5087 24731
rect 5023 24671 5027 24727
rect 5027 24671 5083 24727
rect 5083 24671 5087 24727
rect 5023 24667 5087 24671
rect 5495 24727 5559 24731
rect 5495 24671 5499 24727
rect 5499 24671 5555 24727
rect 5555 24671 5559 24727
rect 5495 24667 5559 24671
rect 5927 24727 5991 24731
rect 5927 24671 5931 24727
rect 5931 24671 5987 24727
rect 5987 24671 5991 24727
rect 5927 24667 5991 24671
rect 6271 24715 6335 24719
rect 6271 24659 6275 24715
rect 6275 24659 6331 24715
rect 6331 24659 6335 24715
rect 6271 24655 6335 24659
rect 6695 24715 6759 24719
rect 6695 24659 6699 24715
rect 6699 24659 6755 24715
rect 6755 24659 6759 24715
rect 6695 24655 6759 24659
rect 5023 24309 5087 24313
rect 5023 24253 5027 24309
rect 5027 24253 5083 24309
rect 5083 24253 5087 24309
rect 5023 24249 5087 24253
rect 5495 24309 5559 24313
rect 5495 24253 5499 24309
rect 5499 24253 5555 24309
rect 5555 24253 5559 24309
rect 5495 24249 5559 24253
rect 5927 24309 5991 24313
rect 5927 24253 5931 24309
rect 5931 24253 5987 24309
rect 5987 24253 5991 24309
rect 5927 24249 5991 24253
rect 6271 24321 6335 24325
rect 6271 24265 6275 24321
rect 6275 24265 6331 24321
rect 6331 24265 6335 24321
rect 6271 24261 6335 24265
rect 6695 24321 6759 24325
rect 6695 24265 6699 24321
rect 6699 24265 6755 24321
rect 6755 24265 6759 24321
rect 6695 24261 6759 24265
rect 5023 23937 5087 23941
rect 5023 23881 5027 23937
rect 5027 23881 5083 23937
rect 5083 23881 5087 23937
rect 5023 23877 5087 23881
rect 5495 23937 5559 23941
rect 5495 23881 5499 23937
rect 5499 23881 5555 23937
rect 5555 23881 5559 23937
rect 5495 23877 5559 23881
rect 5927 23937 5991 23941
rect 5927 23881 5931 23937
rect 5931 23881 5987 23937
rect 5987 23881 5991 23937
rect 5927 23877 5991 23881
rect 6271 23925 6335 23929
rect 6271 23869 6275 23925
rect 6275 23869 6331 23925
rect 6331 23869 6335 23925
rect 6271 23865 6335 23869
rect 6695 23925 6759 23929
rect 6695 23869 6699 23925
rect 6699 23869 6755 23925
rect 6755 23869 6759 23925
rect 6695 23865 6759 23869
rect 5023 23519 5087 23523
rect 5023 23463 5027 23519
rect 5027 23463 5083 23519
rect 5083 23463 5087 23519
rect 5023 23459 5087 23463
rect 5495 23519 5559 23523
rect 5495 23463 5499 23519
rect 5499 23463 5555 23519
rect 5555 23463 5559 23519
rect 5495 23459 5559 23463
rect 5927 23519 5991 23523
rect 5927 23463 5931 23519
rect 5931 23463 5987 23519
rect 5987 23463 5991 23519
rect 5927 23459 5991 23463
rect 6271 23531 6335 23535
rect 6271 23475 6275 23531
rect 6275 23475 6331 23531
rect 6331 23475 6335 23531
rect 6271 23471 6335 23475
rect 6695 23531 6759 23535
rect 6695 23475 6699 23531
rect 6699 23475 6755 23531
rect 6755 23475 6759 23531
rect 6695 23471 6759 23475
rect 5023 23147 5087 23151
rect 5023 23091 5027 23147
rect 5027 23091 5083 23147
rect 5083 23091 5087 23147
rect 5023 23087 5087 23091
rect 5495 23147 5559 23151
rect 5495 23091 5499 23147
rect 5499 23091 5555 23147
rect 5555 23091 5559 23147
rect 5495 23087 5559 23091
rect 5927 23147 5991 23151
rect 5927 23091 5931 23147
rect 5931 23091 5987 23147
rect 5987 23091 5991 23147
rect 5927 23087 5991 23091
rect 6271 23135 6335 23139
rect 6271 23079 6275 23135
rect 6275 23079 6331 23135
rect 6331 23079 6335 23135
rect 6271 23075 6335 23079
rect 6695 23135 6759 23139
rect 6695 23079 6699 23135
rect 6699 23079 6755 23135
rect 6755 23079 6759 23135
rect 6695 23075 6759 23079
rect 5023 22729 5087 22733
rect 5023 22673 5027 22729
rect 5027 22673 5083 22729
rect 5083 22673 5087 22729
rect 5023 22669 5087 22673
rect 5495 22729 5559 22733
rect 5495 22673 5499 22729
rect 5499 22673 5555 22729
rect 5555 22673 5559 22729
rect 5495 22669 5559 22673
rect 5927 22729 5991 22733
rect 5927 22673 5931 22729
rect 5931 22673 5987 22729
rect 5987 22673 5991 22729
rect 5927 22669 5991 22673
rect 6271 22741 6335 22745
rect 6271 22685 6275 22741
rect 6275 22685 6331 22741
rect 6331 22685 6335 22741
rect 6271 22681 6335 22685
rect 6695 22741 6759 22745
rect 6695 22685 6699 22741
rect 6699 22685 6755 22741
rect 6755 22685 6759 22741
rect 6695 22681 6759 22685
rect 5023 22357 5087 22361
rect 5023 22301 5027 22357
rect 5027 22301 5083 22357
rect 5083 22301 5087 22357
rect 5023 22297 5087 22301
rect 5495 22357 5559 22361
rect 5495 22301 5499 22357
rect 5499 22301 5555 22357
rect 5555 22301 5559 22357
rect 5495 22297 5559 22301
rect 5927 22357 5991 22361
rect 5927 22301 5931 22357
rect 5931 22301 5987 22357
rect 5987 22301 5991 22357
rect 5927 22297 5991 22301
rect 6271 22345 6335 22349
rect 6271 22289 6275 22345
rect 6275 22289 6331 22345
rect 6331 22289 6335 22345
rect 6271 22285 6335 22289
rect 6695 22345 6759 22349
rect 6695 22289 6699 22345
rect 6699 22289 6755 22345
rect 6755 22289 6759 22345
rect 6695 22285 6759 22289
rect 5023 21939 5087 21943
rect 5023 21883 5027 21939
rect 5027 21883 5083 21939
rect 5083 21883 5087 21939
rect 5023 21879 5087 21883
rect 5495 21939 5559 21943
rect 5495 21883 5499 21939
rect 5499 21883 5555 21939
rect 5555 21883 5559 21939
rect 5495 21879 5559 21883
rect 5927 21939 5991 21943
rect 5927 21883 5931 21939
rect 5931 21883 5987 21939
rect 5987 21883 5991 21939
rect 5927 21879 5991 21883
rect 6271 21951 6335 21955
rect 6271 21895 6275 21951
rect 6275 21895 6331 21951
rect 6331 21895 6335 21951
rect 6271 21891 6335 21895
rect 6695 21951 6759 21955
rect 6695 21895 6699 21951
rect 6699 21895 6755 21951
rect 6755 21895 6759 21951
rect 6695 21891 6759 21895
rect 5023 21567 5087 21571
rect 5023 21511 5027 21567
rect 5027 21511 5083 21567
rect 5083 21511 5087 21567
rect 5023 21507 5087 21511
rect 5495 21567 5559 21571
rect 5495 21511 5499 21567
rect 5499 21511 5555 21567
rect 5555 21511 5559 21567
rect 5495 21507 5559 21511
rect 5927 21567 5991 21571
rect 5927 21511 5931 21567
rect 5931 21511 5987 21567
rect 5987 21511 5991 21567
rect 5927 21507 5991 21511
rect 6271 21555 6335 21559
rect 6271 21499 6275 21555
rect 6275 21499 6331 21555
rect 6331 21499 6335 21555
rect 6271 21495 6335 21499
rect 6695 21555 6759 21559
rect 6695 21499 6699 21555
rect 6699 21499 6755 21555
rect 6755 21499 6759 21555
rect 6695 21495 6759 21499
rect 5023 21149 5087 21153
rect 5023 21093 5027 21149
rect 5027 21093 5083 21149
rect 5083 21093 5087 21149
rect 5023 21089 5087 21093
rect 5495 21149 5559 21153
rect 5495 21093 5499 21149
rect 5499 21093 5555 21149
rect 5555 21093 5559 21149
rect 5495 21089 5559 21093
rect 5927 21149 5991 21153
rect 5927 21093 5931 21149
rect 5931 21093 5987 21149
rect 5987 21093 5991 21149
rect 5927 21089 5991 21093
rect 6271 21161 6335 21165
rect 6271 21105 6275 21161
rect 6275 21105 6331 21161
rect 6331 21105 6335 21161
rect 6271 21101 6335 21105
rect 6695 21161 6759 21165
rect 6695 21105 6699 21161
rect 6699 21105 6755 21161
rect 6755 21105 6759 21161
rect 6695 21101 6759 21105
rect 5023 20777 5087 20781
rect 5023 20721 5027 20777
rect 5027 20721 5083 20777
rect 5083 20721 5087 20777
rect 5023 20717 5087 20721
rect 5495 20777 5559 20781
rect 5495 20721 5499 20777
rect 5499 20721 5555 20777
rect 5555 20721 5559 20777
rect 5495 20717 5559 20721
rect 5927 20777 5991 20781
rect 5927 20721 5931 20777
rect 5931 20721 5987 20777
rect 5987 20721 5991 20777
rect 5927 20717 5991 20721
rect 6271 20765 6335 20769
rect 6271 20709 6275 20765
rect 6275 20709 6331 20765
rect 6331 20709 6335 20765
rect 6271 20705 6335 20709
rect 6695 20765 6759 20769
rect 6695 20709 6699 20765
rect 6699 20709 6755 20765
rect 6755 20709 6759 20765
rect 6695 20705 6759 20709
rect 5023 20359 5087 20363
rect 5023 20303 5027 20359
rect 5027 20303 5083 20359
rect 5083 20303 5087 20359
rect 5023 20299 5087 20303
rect 5495 20359 5559 20363
rect 5495 20303 5499 20359
rect 5499 20303 5555 20359
rect 5555 20303 5559 20359
rect 5495 20299 5559 20303
rect 5927 20359 5991 20363
rect 5927 20303 5931 20359
rect 5931 20303 5987 20359
rect 5987 20303 5991 20359
rect 5927 20299 5991 20303
rect 6271 20371 6335 20375
rect 6271 20315 6275 20371
rect 6275 20315 6331 20371
rect 6331 20315 6335 20371
rect 6271 20311 6335 20315
rect 6695 20371 6759 20375
rect 6695 20315 6699 20371
rect 6699 20315 6755 20371
rect 6755 20315 6759 20371
rect 6695 20311 6759 20315
rect 5023 19987 5087 19991
rect 5023 19931 5027 19987
rect 5027 19931 5083 19987
rect 5083 19931 5087 19987
rect 5023 19927 5087 19931
rect 5495 19987 5559 19991
rect 5495 19931 5499 19987
rect 5499 19931 5555 19987
rect 5555 19931 5559 19987
rect 5495 19927 5559 19931
rect 5927 19987 5991 19991
rect 5927 19931 5931 19987
rect 5931 19931 5987 19987
rect 5987 19931 5991 19987
rect 5927 19927 5991 19931
rect 6271 19975 6335 19979
rect 6271 19919 6275 19975
rect 6275 19919 6331 19975
rect 6331 19919 6335 19975
rect 6271 19915 6335 19919
rect 6695 19975 6759 19979
rect 6695 19919 6699 19975
rect 6699 19919 6755 19975
rect 6755 19919 6759 19975
rect 6695 19915 6759 19919
rect 5023 19569 5087 19573
rect 5023 19513 5027 19569
rect 5027 19513 5083 19569
rect 5083 19513 5087 19569
rect 5023 19509 5087 19513
rect 5495 19569 5559 19573
rect 5495 19513 5499 19569
rect 5499 19513 5555 19569
rect 5555 19513 5559 19569
rect 5495 19509 5559 19513
rect 5927 19569 5991 19573
rect 5927 19513 5931 19569
rect 5931 19513 5987 19569
rect 5987 19513 5991 19569
rect 5927 19509 5991 19513
rect 6271 19581 6335 19585
rect 6271 19525 6275 19581
rect 6275 19525 6331 19581
rect 6331 19525 6335 19581
rect 6271 19521 6335 19525
rect 6695 19581 6759 19585
rect 6695 19525 6699 19581
rect 6699 19525 6755 19581
rect 6755 19525 6759 19581
rect 6695 19521 6759 19525
rect 5023 19197 5087 19201
rect 5023 19141 5027 19197
rect 5027 19141 5083 19197
rect 5083 19141 5087 19197
rect 5023 19137 5087 19141
rect 5495 19197 5559 19201
rect 5495 19141 5499 19197
rect 5499 19141 5555 19197
rect 5555 19141 5559 19197
rect 5495 19137 5559 19141
rect 5927 19197 5991 19201
rect 5927 19141 5931 19197
rect 5931 19141 5987 19197
rect 5987 19141 5991 19197
rect 5927 19137 5991 19141
rect 6271 19185 6335 19189
rect 6271 19129 6275 19185
rect 6275 19129 6331 19185
rect 6331 19129 6335 19185
rect 6271 19125 6335 19129
rect 6695 19185 6759 19189
rect 6695 19129 6699 19185
rect 6699 19129 6755 19185
rect 6755 19129 6759 19185
rect 6695 19125 6759 19129
rect 5023 18779 5087 18783
rect 5023 18723 5027 18779
rect 5027 18723 5083 18779
rect 5083 18723 5087 18779
rect 5023 18719 5087 18723
rect 5495 18779 5559 18783
rect 5495 18723 5499 18779
rect 5499 18723 5555 18779
rect 5555 18723 5559 18779
rect 5495 18719 5559 18723
rect 5927 18779 5991 18783
rect 5927 18723 5931 18779
rect 5931 18723 5987 18779
rect 5987 18723 5991 18779
rect 5927 18719 5991 18723
rect 6271 18791 6335 18795
rect 6271 18735 6275 18791
rect 6275 18735 6331 18791
rect 6331 18735 6335 18791
rect 6271 18731 6335 18735
rect 6695 18791 6759 18795
rect 6695 18735 6699 18791
rect 6699 18735 6755 18791
rect 6755 18735 6759 18791
rect 6695 18731 6759 18735
rect 5023 18407 5087 18411
rect 5023 18351 5027 18407
rect 5027 18351 5083 18407
rect 5083 18351 5087 18407
rect 5023 18347 5087 18351
rect 5495 18407 5559 18411
rect 5495 18351 5499 18407
rect 5499 18351 5555 18407
rect 5555 18351 5559 18407
rect 5495 18347 5559 18351
rect 5927 18407 5991 18411
rect 5927 18351 5931 18407
rect 5931 18351 5987 18407
rect 5987 18351 5991 18407
rect 5927 18347 5991 18351
rect 6271 18395 6335 18399
rect 6271 18339 6275 18395
rect 6275 18339 6331 18395
rect 6331 18339 6335 18395
rect 6271 18335 6335 18339
rect 6695 18395 6759 18399
rect 6695 18339 6699 18395
rect 6699 18339 6755 18395
rect 6755 18339 6759 18395
rect 6695 18335 6759 18339
rect 5023 17989 5087 17993
rect 5023 17933 5027 17989
rect 5027 17933 5083 17989
rect 5083 17933 5087 17989
rect 5023 17929 5087 17933
rect 5495 17989 5559 17993
rect 5495 17933 5499 17989
rect 5499 17933 5555 17989
rect 5555 17933 5559 17989
rect 5495 17929 5559 17933
rect 5927 17989 5991 17993
rect 5927 17933 5931 17989
rect 5931 17933 5987 17989
rect 5987 17933 5991 17989
rect 5927 17929 5991 17933
rect 6271 18001 6335 18005
rect 6271 17945 6275 18001
rect 6275 17945 6331 18001
rect 6331 17945 6335 18001
rect 6271 17941 6335 17945
rect 6695 18001 6759 18005
rect 6695 17945 6699 18001
rect 6699 17945 6755 18001
rect 6755 17945 6759 18001
rect 6695 17941 6759 17945
rect 5023 17617 5087 17621
rect 5023 17561 5027 17617
rect 5027 17561 5083 17617
rect 5083 17561 5087 17617
rect 5023 17557 5087 17561
rect 5495 17617 5559 17621
rect 5495 17561 5499 17617
rect 5499 17561 5555 17617
rect 5555 17561 5559 17617
rect 5495 17557 5559 17561
rect 5927 17617 5991 17621
rect 5927 17561 5931 17617
rect 5931 17561 5987 17617
rect 5987 17561 5991 17617
rect 5927 17557 5991 17561
rect 6271 17605 6335 17609
rect 6271 17549 6275 17605
rect 6275 17549 6331 17605
rect 6331 17549 6335 17605
rect 6271 17545 6335 17549
rect 6695 17605 6759 17609
rect 6695 17549 6699 17605
rect 6699 17549 6755 17605
rect 6755 17549 6759 17605
rect 6695 17545 6759 17549
rect 5023 17199 5087 17203
rect 5023 17143 5027 17199
rect 5027 17143 5083 17199
rect 5083 17143 5087 17199
rect 5023 17139 5087 17143
rect 5495 17199 5559 17203
rect 5495 17143 5499 17199
rect 5499 17143 5555 17199
rect 5555 17143 5559 17199
rect 5495 17139 5559 17143
rect 5927 17199 5991 17203
rect 5927 17143 5931 17199
rect 5931 17143 5987 17199
rect 5987 17143 5991 17199
rect 5927 17139 5991 17143
rect 6271 17211 6335 17215
rect 6271 17155 6275 17211
rect 6275 17155 6331 17211
rect 6331 17155 6335 17211
rect 6271 17151 6335 17155
rect 6695 17211 6759 17215
rect 6695 17155 6699 17211
rect 6699 17155 6755 17211
rect 6755 17155 6759 17211
rect 6695 17151 6759 17155
rect 5023 16827 5087 16831
rect 5023 16771 5027 16827
rect 5027 16771 5083 16827
rect 5083 16771 5087 16827
rect 5023 16767 5087 16771
rect 5495 16827 5559 16831
rect 5495 16771 5499 16827
rect 5499 16771 5555 16827
rect 5555 16771 5559 16827
rect 5495 16767 5559 16771
rect 5927 16827 5991 16831
rect 5927 16771 5931 16827
rect 5931 16771 5987 16827
rect 5987 16771 5991 16827
rect 5927 16767 5991 16771
rect 6271 16815 6335 16819
rect 6271 16759 6275 16815
rect 6275 16759 6331 16815
rect 6331 16759 6335 16815
rect 6271 16755 6335 16759
rect 6695 16815 6759 16819
rect 6695 16759 6699 16815
rect 6699 16759 6755 16815
rect 6755 16759 6759 16815
rect 6695 16755 6759 16759
rect 5023 16409 5087 16413
rect 5023 16353 5027 16409
rect 5027 16353 5083 16409
rect 5083 16353 5087 16409
rect 5023 16349 5087 16353
rect 5495 16409 5559 16413
rect 5495 16353 5499 16409
rect 5499 16353 5555 16409
rect 5555 16353 5559 16409
rect 5495 16349 5559 16353
rect 5927 16409 5991 16413
rect 5927 16353 5931 16409
rect 5931 16353 5987 16409
rect 5987 16353 5991 16409
rect 5927 16349 5991 16353
rect 6271 16421 6335 16425
rect 6271 16365 6275 16421
rect 6275 16365 6331 16421
rect 6331 16365 6335 16421
rect 6271 16361 6335 16365
rect 6695 16421 6759 16425
rect 6695 16365 6699 16421
rect 6699 16365 6755 16421
rect 6755 16365 6759 16421
rect 6695 16361 6759 16365
rect 5023 16037 5087 16041
rect 5023 15981 5027 16037
rect 5027 15981 5083 16037
rect 5083 15981 5087 16037
rect 5023 15977 5087 15981
rect 5495 16037 5559 16041
rect 5495 15981 5499 16037
rect 5499 15981 5555 16037
rect 5555 15981 5559 16037
rect 5495 15977 5559 15981
rect 5927 16037 5991 16041
rect 5927 15981 5931 16037
rect 5931 15981 5987 16037
rect 5987 15981 5991 16037
rect 5927 15977 5991 15981
rect 6271 16025 6335 16029
rect 6271 15969 6275 16025
rect 6275 15969 6331 16025
rect 6331 15969 6335 16025
rect 6271 15965 6335 15969
rect 6695 16025 6759 16029
rect 6695 15969 6699 16025
rect 6699 15969 6755 16025
rect 6755 15969 6759 16025
rect 6695 15965 6759 15969
rect 5023 15619 5087 15623
rect 5023 15563 5027 15619
rect 5027 15563 5083 15619
rect 5083 15563 5087 15619
rect 5023 15559 5087 15563
rect 5495 15619 5559 15623
rect 5495 15563 5499 15619
rect 5499 15563 5555 15619
rect 5555 15563 5559 15619
rect 5495 15559 5559 15563
rect 5927 15619 5991 15623
rect 5927 15563 5931 15619
rect 5931 15563 5987 15619
rect 5987 15563 5991 15619
rect 5927 15559 5991 15563
rect 6271 15631 6335 15635
rect 6271 15575 6275 15631
rect 6275 15575 6331 15631
rect 6331 15575 6335 15631
rect 6271 15571 6335 15575
rect 6695 15631 6759 15635
rect 6695 15575 6699 15631
rect 6699 15575 6755 15631
rect 6755 15575 6759 15631
rect 6695 15571 6759 15575
rect 5023 15247 5087 15251
rect 5023 15191 5027 15247
rect 5027 15191 5083 15247
rect 5083 15191 5087 15247
rect 5023 15187 5087 15191
rect 5495 15247 5559 15251
rect 5495 15191 5499 15247
rect 5499 15191 5555 15247
rect 5555 15191 5559 15247
rect 5495 15187 5559 15191
rect 5927 15247 5991 15251
rect 5927 15191 5931 15247
rect 5931 15191 5987 15247
rect 5987 15191 5991 15247
rect 5927 15187 5991 15191
rect 6271 15235 6335 15239
rect 6271 15179 6275 15235
rect 6275 15179 6331 15235
rect 6331 15179 6335 15235
rect 6271 15175 6335 15179
rect 6695 15235 6759 15239
rect 6695 15179 6699 15235
rect 6699 15179 6755 15235
rect 6755 15179 6759 15235
rect 6695 15175 6759 15179
rect 5023 14829 5087 14833
rect 5023 14773 5027 14829
rect 5027 14773 5083 14829
rect 5083 14773 5087 14829
rect 5023 14769 5087 14773
rect 5495 14829 5559 14833
rect 5495 14773 5499 14829
rect 5499 14773 5555 14829
rect 5555 14773 5559 14829
rect 5495 14769 5559 14773
rect 5927 14829 5991 14833
rect 5927 14773 5931 14829
rect 5931 14773 5987 14829
rect 5987 14773 5991 14829
rect 5927 14769 5991 14773
rect 6271 14841 6335 14845
rect 6271 14785 6275 14841
rect 6275 14785 6331 14841
rect 6331 14785 6335 14841
rect 6271 14781 6335 14785
rect 6695 14841 6759 14845
rect 6695 14785 6699 14841
rect 6699 14785 6755 14841
rect 6755 14785 6759 14841
rect 6695 14781 6759 14785
rect 5023 14457 5087 14461
rect 5023 14401 5027 14457
rect 5027 14401 5083 14457
rect 5083 14401 5087 14457
rect 5023 14397 5087 14401
rect 5495 14457 5559 14461
rect 5495 14401 5499 14457
rect 5499 14401 5555 14457
rect 5555 14401 5559 14457
rect 5495 14397 5559 14401
rect 5927 14457 5991 14461
rect 5927 14401 5931 14457
rect 5931 14401 5987 14457
rect 5987 14401 5991 14457
rect 5927 14397 5991 14401
rect 6271 14445 6335 14449
rect 6271 14389 6275 14445
rect 6275 14389 6331 14445
rect 6331 14389 6335 14445
rect 6271 14385 6335 14389
rect 6695 14445 6759 14449
rect 6695 14389 6699 14445
rect 6699 14389 6755 14445
rect 6755 14389 6759 14445
rect 6695 14385 6759 14389
rect 5023 14039 5087 14043
rect 5023 13983 5027 14039
rect 5027 13983 5083 14039
rect 5083 13983 5087 14039
rect 5023 13979 5087 13983
rect 5495 14039 5559 14043
rect 5495 13983 5499 14039
rect 5499 13983 5555 14039
rect 5555 13983 5559 14039
rect 5495 13979 5559 13983
rect 5927 14039 5991 14043
rect 5927 13983 5931 14039
rect 5931 13983 5987 14039
rect 5987 13983 5991 14039
rect 5927 13979 5991 13983
rect 6271 14051 6335 14055
rect 6271 13995 6275 14051
rect 6275 13995 6331 14051
rect 6331 13995 6335 14051
rect 6271 13991 6335 13995
rect 6695 14051 6759 14055
rect 6695 13995 6699 14051
rect 6699 13995 6755 14051
rect 6755 13995 6759 14051
rect 6695 13991 6759 13995
rect 5023 13667 5087 13671
rect 5023 13611 5027 13667
rect 5027 13611 5083 13667
rect 5083 13611 5087 13667
rect 5023 13607 5087 13611
rect 5495 13667 5559 13671
rect 5495 13611 5499 13667
rect 5499 13611 5555 13667
rect 5555 13611 5559 13667
rect 5495 13607 5559 13611
rect 5927 13667 5991 13671
rect 5927 13611 5931 13667
rect 5931 13611 5987 13667
rect 5987 13611 5991 13667
rect 5927 13607 5991 13611
rect 6271 13655 6335 13659
rect 6271 13599 6275 13655
rect 6275 13599 6331 13655
rect 6331 13599 6335 13655
rect 6271 13595 6335 13599
rect 6695 13655 6759 13659
rect 6695 13599 6699 13655
rect 6699 13599 6755 13655
rect 6755 13599 6759 13655
rect 6695 13595 6759 13599
rect 5023 13249 5087 13253
rect 5023 13193 5027 13249
rect 5027 13193 5083 13249
rect 5083 13193 5087 13249
rect 5023 13189 5087 13193
rect 5495 13249 5559 13253
rect 5495 13193 5499 13249
rect 5499 13193 5555 13249
rect 5555 13193 5559 13249
rect 5495 13189 5559 13193
rect 5927 13249 5991 13253
rect 5927 13193 5931 13249
rect 5931 13193 5987 13249
rect 5987 13193 5991 13249
rect 5927 13189 5991 13193
rect 6271 13261 6335 13265
rect 6271 13205 6275 13261
rect 6275 13205 6331 13261
rect 6331 13205 6335 13261
rect 6271 13201 6335 13205
rect 6695 13261 6759 13265
rect 6695 13205 6699 13261
rect 6699 13205 6755 13261
rect 6755 13205 6759 13261
rect 6695 13201 6759 13205
rect 5023 12877 5087 12881
rect 5023 12821 5027 12877
rect 5027 12821 5083 12877
rect 5083 12821 5087 12877
rect 5023 12817 5087 12821
rect 5495 12877 5559 12881
rect 5495 12821 5499 12877
rect 5499 12821 5555 12877
rect 5555 12821 5559 12877
rect 5495 12817 5559 12821
rect 5927 12877 5991 12881
rect 5927 12821 5931 12877
rect 5931 12821 5987 12877
rect 5987 12821 5991 12877
rect 5927 12817 5991 12821
rect 6271 12865 6335 12869
rect 6271 12809 6275 12865
rect 6275 12809 6331 12865
rect 6331 12809 6335 12865
rect 6271 12805 6335 12809
rect 6695 12865 6759 12869
rect 6695 12809 6699 12865
rect 6699 12809 6755 12865
rect 6755 12809 6759 12865
rect 6695 12805 6759 12809
rect 5023 12459 5087 12463
rect 5023 12403 5027 12459
rect 5027 12403 5083 12459
rect 5083 12403 5087 12459
rect 5023 12399 5087 12403
rect 5495 12459 5559 12463
rect 5495 12403 5499 12459
rect 5499 12403 5555 12459
rect 5555 12403 5559 12459
rect 5495 12399 5559 12403
rect 5927 12459 5991 12463
rect 5927 12403 5931 12459
rect 5931 12403 5987 12459
rect 5987 12403 5991 12459
rect 5927 12399 5991 12403
rect 6271 12471 6335 12475
rect 6271 12415 6275 12471
rect 6275 12415 6331 12471
rect 6331 12415 6335 12471
rect 6271 12411 6335 12415
rect 6695 12471 6759 12475
rect 6695 12415 6699 12471
rect 6699 12415 6755 12471
rect 6755 12415 6759 12471
rect 6695 12411 6759 12415
rect 5023 12087 5087 12091
rect 5023 12031 5027 12087
rect 5027 12031 5083 12087
rect 5083 12031 5087 12087
rect 5023 12027 5087 12031
rect 5495 12087 5559 12091
rect 5495 12031 5499 12087
rect 5499 12031 5555 12087
rect 5555 12031 5559 12087
rect 5495 12027 5559 12031
rect 5927 12087 5991 12091
rect 5927 12031 5931 12087
rect 5931 12031 5987 12087
rect 5987 12031 5991 12087
rect 5927 12027 5991 12031
rect 6271 12075 6335 12079
rect 6271 12019 6275 12075
rect 6275 12019 6331 12075
rect 6331 12019 6335 12075
rect 6271 12015 6335 12019
rect 6695 12075 6759 12079
rect 6695 12019 6699 12075
rect 6699 12019 6755 12075
rect 6755 12019 6759 12075
rect 6695 12015 6759 12019
rect 5023 11669 5087 11673
rect 5023 11613 5027 11669
rect 5027 11613 5083 11669
rect 5083 11613 5087 11669
rect 5023 11609 5087 11613
rect 5495 11669 5559 11673
rect 5495 11613 5499 11669
rect 5499 11613 5555 11669
rect 5555 11613 5559 11669
rect 5495 11609 5559 11613
rect 5927 11669 5991 11673
rect 5927 11613 5931 11669
rect 5931 11613 5987 11669
rect 5987 11613 5991 11669
rect 5927 11609 5991 11613
rect 6271 11681 6335 11685
rect 6271 11625 6275 11681
rect 6275 11625 6331 11681
rect 6331 11625 6335 11681
rect 6271 11621 6335 11625
rect 6695 11681 6759 11685
rect 6695 11625 6699 11681
rect 6699 11625 6755 11681
rect 6755 11625 6759 11681
rect 6695 11621 6759 11625
rect 5023 11297 5087 11301
rect 5023 11241 5027 11297
rect 5027 11241 5083 11297
rect 5083 11241 5087 11297
rect 5023 11237 5087 11241
rect 5495 11297 5559 11301
rect 5495 11241 5499 11297
rect 5499 11241 5555 11297
rect 5555 11241 5559 11297
rect 5495 11237 5559 11241
rect 5927 11297 5991 11301
rect 5927 11241 5931 11297
rect 5931 11241 5987 11297
rect 5987 11241 5991 11297
rect 5927 11237 5991 11241
rect 6271 11285 6335 11289
rect 6271 11229 6275 11285
rect 6275 11229 6331 11285
rect 6331 11229 6335 11285
rect 6271 11225 6335 11229
rect 6695 11285 6759 11289
rect 6695 11229 6699 11285
rect 6699 11229 6755 11285
rect 6755 11229 6759 11285
rect 6695 11225 6759 11229
rect 5023 10879 5087 10883
rect 5023 10823 5027 10879
rect 5027 10823 5083 10879
rect 5083 10823 5087 10879
rect 5023 10819 5087 10823
rect 5495 10879 5559 10883
rect 5495 10823 5499 10879
rect 5499 10823 5555 10879
rect 5555 10823 5559 10879
rect 5495 10819 5559 10823
rect 5927 10879 5991 10883
rect 5927 10823 5931 10879
rect 5931 10823 5987 10879
rect 5987 10823 5991 10879
rect 5927 10819 5991 10823
rect 6271 10891 6335 10895
rect 6271 10835 6275 10891
rect 6275 10835 6331 10891
rect 6331 10835 6335 10891
rect 6271 10831 6335 10835
rect 6695 10891 6759 10895
rect 6695 10835 6699 10891
rect 6699 10835 6755 10891
rect 6755 10835 6759 10891
rect 6695 10831 6759 10835
rect 5023 10507 5087 10511
rect 5023 10451 5027 10507
rect 5027 10451 5083 10507
rect 5083 10451 5087 10507
rect 5023 10447 5087 10451
rect 5495 10507 5559 10511
rect 5495 10451 5499 10507
rect 5499 10451 5555 10507
rect 5555 10451 5559 10507
rect 5495 10447 5559 10451
rect 5927 10507 5991 10511
rect 5927 10451 5931 10507
rect 5931 10451 5987 10507
rect 5987 10451 5991 10507
rect 5927 10447 5991 10451
rect 6271 10495 6335 10499
rect 6271 10439 6275 10495
rect 6275 10439 6331 10495
rect 6331 10439 6335 10495
rect 6271 10435 6335 10439
rect 6695 10495 6759 10499
rect 6695 10439 6699 10495
rect 6699 10439 6755 10495
rect 6755 10439 6759 10495
rect 6695 10435 6759 10439
rect 5023 10089 5087 10093
rect 5023 10033 5027 10089
rect 5027 10033 5083 10089
rect 5083 10033 5087 10089
rect 5023 10029 5087 10033
rect 5495 10089 5559 10093
rect 5495 10033 5499 10089
rect 5499 10033 5555 10089
rect 5555 10033 5559 10089
rect 5495 10029 5559 10033
rect 5927 10089 5991 10093
rect 5927 10033 5931 10089
rect 5931 10033 5987 10089
rect 5987 10033 5991 10089
rect 5927 10029 5991 10033
rect 6271 10101 6335 10105
rect 6271 10045 6275 10101
rect 6275 10045 6331 10101
rect 6331 10045 6335 10101
rect 6271 10041 6335 10045
rect 6695 10101 6759 10105
rect 6695 10045 6699 10101
rect 6699 10045 6755 10101
rect 6755 10045 6759 10101
rect 6695 10041 6759 10045
rect 5023 9717 5087 9721
rect 5023 9661 5027 9717
rect 5027 9661 5083 9717
rect 5083 9661 5087 9717
rect 5023 9657 5087 9661
rect 5495 9717 5559 9721
rect 5495 9661 5499 9717
rect 5499 9661 5555 9717
rect 5555 9661 5559 9717
rect 5495 9657 5559 9661
rect 5927 9717 5991 9721
rect 5927 9661 5931 9717
rect 5931 9661 5987 9717
rect 5987 9661 5991 9717
rect 5927 9657 5991 9661
rect 6271 9705 6335 9709
rect 6271 9649 6275 9705
rect 6275 9649 6331 9705
rect 6331 9649 6335 9705
rect 6271 9645 6335 9649
rect 6695 9705 6759 9709
rect 6695 9649 6699 9705
rect 6699 9649 6755 9705
rect 6755 9649 6759 9705
rect 6695 9645 6759 9649
rect 5023 9299 5087 9303
rect 5023 9243 5027 9299
rect 5027 9243 5083 9299
rect 5083 9243 5087 9299
rect 5023 9239 5087 9243
rect 5495 9299 5559 9303
rect 5495 9243 5499 9299
rect 5499 9243 5555 9299
rect 5555 9243 5559 9299
rect 5495 9239 5559 9243
rect 5927 9299 5991 9303
rect 5927 9243 5931 9299
rect 5931 9243 5987 9299
rect 5987 9243 5991 9299
rect 5927 9239 5991 9243
rect 6271 9311 6335 9315
rect 6271 9255 6275 9311
rect 6275 9255 6331 9311
rect 6331 9255 6335 9311
rect 6271 9251 6335 9255
rect 6695 9311 6759 9315
rect 6695 9255 6699 9311
rect 6699 9255 6755 9311
rect 6755 9255 6759 9311
rect 6695 9251 6759 9255
rect 5023 8927 5087 8931
rect 5023 8871 5027 8927
rect 5027 8871 5083 8927
rect 5083 8871 5087 8927
rect 5023 8867 5087 8871
rect 5495 8927 5559 8931
rect 5495 8871 5499 8927
rect 5499 8871 5555 8927
rect 5555 8871 5559 8927
rect 5495 8867 5559 8871
rect 5927 8927 5991 8931
rect 5927 8871 5931 8927
rect 5931 8871 5987 8927
rect 5987 8871 5991 8927
rect 5927 8867 5991 8871
rect 6271 8915 6335 8919
rect 6271 8859 6275 8915
rect 6275 8859 6331 8915
rect 6331 8859 6335 8915
rect 6271 8855 6335 8859
rect 6695 8915 6759 8919
rect 6695 8859 6699 8915
rect 6699 8859 6755 8915
rect 6755 8859 6759 8915
rect 6695 8855 6759 8859
rect 5023 8509 5087 8513
rect 5023 8453 5027 8509
rect 5027 8453 5083 8509
rect 5083 8453 5087 8509
rect 5023 8449 5087 8453
rect 5495 8509 5559 8513
rect 5495 8453 5499 8509
rect 5499 8453 5555 8509
rect 5555 8453 5559 8509
rect 5495 8449 5559 8453
rect 5927 8509 5991 8513
rect 5927 8453 5931 8509
rect 5931 8453 5987 8509
rect 5987 8453 5991 8509
rect 5927 8449 5991 8453
rect 6271 8521 6335 8525
rect 6271 8465 6275 8521
rect 6275 8465 6331 8521
rect 6331 8465 6335 8521
rect 6271 8461 6335 8465
rect 6695 8521 6759 8525
rect 6695 8465 6699 8521
rect 6699 8465 6755 8521
rect 6755 8465 6759 8521
rect 6695 8461 6759 8465
rect 5023 8137 5087 8141
rect 5023 8081 5027 8137
rect 5027 8081 5083 8137
rect 5083 8081 5087 8137
rect 5023 8077 5087 8081
rect 5495 8137 5559 8141
rect 5495 8081 5499 8137
rect 5499 8081 5555 8137
rect 5555 8081 5559 8137
rect 5495 8077 5559 8081
rect 5927 8137 5991 8141
rect 5927 8081 5931 8137
rect 5931 8081 5987 8137
rect 5987 8081 5991 8137
rect 5927 8077 5991 8081
rect 6271 8125 6335 8129
rect 6271 8069 6275 8125
rect 6275 8069 6331 8125
rect 6331 8069 6335 8125
rect 6271 8065 6335 8069
rect 6695 8125 6759 8129
rect 6695 8069 6699 8125
rect 6699 8069 6755 8125
rect 6755 8069 6759 8125
rect 6695 8065 6759 8069
rect 5023 7719 5087 7723
rect 5023 7663 5027 7719
rect 5027 7663 5083 7719
rect 5083 7663 5087 7719
rect 5023 7659 5087 7663
rect 5495 7719 5559 7723
rect 5495 7663 5499 7719
rect 5499 7663 5555 7719
rect 5555 7663 5559 7719
rect 5495 7659 5559 7663
rect 5927 7719 5991 7723
rect 5927 7663 5931 7719
rect 5931 7663 5987 7719
rect 5987 7663 5991 7719
rect 5927 7659 5991 7663
rect 6271 7731 6335 7735
rect 6271 7675 6275 7731
rect 6275 7675 6331 7731
rect 6331 7675 6335 7731
rect 6271 7671 6335 7675
rect 6695 7731 6759 7735
rect 6695 7675 6699 7731
rect 6699 7675 6755 7731
rect 6755 7675 6759 7731
rect 6695 7671 6759 7675
rect 5023 7347 5087 7351
rect 5023 7291 5027 7347
rect 5027 7291 5083 7347
rect 5083 7291 5087 7347
rect 5023 7287 5087 7291
rect 5495 7347 5559 7351
rect 5495 7291 5499 7347
rect 5499 7291 5555 7347
rect 5555 7291 5559 7347
rect 5495 7287 5559 7291
rect 5927 7347 5991 7351
rect 5927 7291 5931 7347
rect 5931 7291 5987 7347
rect 5987 7291 5991 7347
rect 5927 7287 5991 7291
rect 6271 7335 6335 7339
rect 6271 7279 6275 7335
rect 6275 7279 6331 7335
rect 6331 7279 6335 7335
rect 6271 7275 6335 7279
rect 6695 7335 6759 7339
rect 6695 7279 6699 7335
rect 6699 7279 6755 7335
rect 6755 7279 6759 7335
rect 6695 7275 6759 7279
rect 5023 6929 5087 6933
rect 5023 6873 5027 6929
rect 5027 6873 5083 6929
rect 5083 6873 5087 6929
rect 5023 6869 5087 6873
rect 5495 6929 5559 6933
rect 5495 6873 5499 6929
rect 5499 6873 5555 6929
rect 5555 6873 5559 6929
rect 5495 6869 5559 6873
rect 5927 6929 5991 6933
rect 5927 6873 5931 6929
rect 5931 6873 5987 6929
rect 5987 6873 5991 6929
rect 5927 6869 5991 6873
rect 6271 6941 6335 6945
rect 6271 6885 6275 6941
rect 6275 6885 6331 6941
rect 6331 6885 6335 6941
rect 6271 6881 6335 6885
rect 6695 6941 6759 6945
rect 6695 6885 6699 6941
rect 6699 6885 6755 6941
rect 6755 6885 6759 6941
rect 6695 6881 6759 6885
rect 5023 6557 5087 6561
rect 5023 6501 5027 6557
rect 5027 6501 5083 6557
rect 5083 6501 5087 6557
rect 5023 6497 5087 6501
rect 5495 6557 5559 6561
rect 5495 6501 5499 6557
rect 5499 6501 5555 6557
rect 5555 6501 5559 6557
rect 5495 6497 5559 6501
rect 5927 6557 5991 6561
rect 5927 6501 5931 6557
rect 5931 6501 5987 6557
rect 5987 6501 5991 6557
rect 5927 6497 5991 6501
rect 6271 6545 6335 6549
rect 6271 6489 6275 6545
rect 6275 6489 6331 6545
rect 6331 6489 6335 6545
rect 6271 6485 6335 6489
rect 6695 6545 6759 6549
rect 6695 6489 6699 6545
rect 6699 6489 6755 6545
rect 6755 6489 6759 6545
rect 6695 6485 6759 6489
rect 5023 6139 5087 6143
rect 5023 6083 5027 6139
rect 5027 6083 5083 6139
rect 5083 6083 5087 6139
rect 5023 6079 5087 6083
rect 5495 6139 5559 6143
rect 5495 6083 5499 6139
rect 5499 6083 5555 6139
rect 5555 6083 5559 6139
rect 5495 6079 5559 6083
rect 5927 6139 5991 6143
rect 5927 6083 5931 6139
rect 5931 6083 5987 6139
rect 5987 6083 5991 6139
rect 5927 6079 5991 6083
rect 6271 6151 6335 6155
rect 6271 6095 6275 6151
rect 6275 6095 6331 6151
rect 6331 6095 6335 6151
rect 6271 6091 6335 6095
rect 6695 6151 6759 6155
rect 6695 6095 6699 6151
rect 6699 6095 6755 6151
rect 6755 6095 6759 6151
rect 6695 6091 6759 6095
rect 5023 5767 5087 5771
rect 5023 5711 5027 5767
rect 5027 5711 5083 5767
rect 5083 5711 5087 5767
rect 5023 5707 5087 5711
rect 5495 5767 5559 5771
rect 5495 5711 5499 5767
rect 5499 5711 5555 5767
rect 5555 5711 5559 5767
rect 5495 5707 5559 5711
rect 5927 5767 5991 5771
rect 5927 5711 5931 5767
rect 5931 5711 5987 5767
rect 5987 5711 5991 5767
rect 5927 5707 5991 5711
rect 6271 5755 6335 5759
rect 6271 5699 6275 5755
rect 6275 5699 6331 5755
rect 6331 5699 6335 5755
rect 6271 5695 6335 5699
rect 6695 5755 6759 5759
rect 6695 5699 6699 5755
rect 6699 5699 6755 5755
rect 6755 5699 6759 5755
rect 6695 5695 6759 5699
rect 5023 5349 5087 5353
rect 5023 5293 5027 5349
rect 5027 5293 5083 5349
rect 5083 5293 5087 5349
rect 5023 5289 5087 5293
rect 5495 5349 5559 5353
rect 5495 5293 5499 5349
rect 5499 5293 5555 5349
rect 5555 5293 5559 5349
rect 5495 5289 5559 5293
rect 5927 5349 5991 5353
rect 5927 5293 5931 5349
rect 5931 5293 5987 5349
rect 5987 5293 5991 5349
rect 5927 5289 5991 5293
rect 6271 5361 6335 5365
rect 6271 5305 6275 5361
rect 6275 5305 6331 5361
rect 6331 5305 6335 5361
rect 6271 5301 6335 5305
rect 6695 5361 6759 5365
rect 6695 5305 6699 5361
rect 6699 5305 6755 5361
rect 6755 5305 6759 5361
rect 6695 5301 6759 5305
rect 5023 4977 5087 4981
rect 5023 4921 5027 4977
rect 5027 4921 5083 4977
rect 5083 4921 5087 4977
rect 5023 4917 5087 4921
rect 5495 4977 5559 4981
rect 5495 4921 5499 4977
rect 5499 4921 5555 4977
rect 5555 4921 5559 4977
rect 5495 4917 5559 4921
rect 5927 4977 5991 4981
rect 5927 4921 5931 4977
rect 5931 4921 5987 4977
rect 5987 4921 5991 4977
rect 5927 4917 5991 4921
rect 6271 4965 6335 4969
rect 6271 4909 6275 4965
rect 6275 4909 6331 4965
rect 6331 4909 6335 4965
rect 6271 4905 6335 4909
rect 6695 4965 6759 4969
rect 6695 4909 6699 4965
rect 6699 4909 6755 4965
rect 6755 4909 6759 4965
rect 6695 4905 6759 4909
rect 5023 4559 5087 4563
rect 5023 4503 5027 4559
rect 5027 4503 5083 4559
rect 5083 4503 5087 4559
rect 5023 4499 5087 4503
rect 5495 4559 5559 4563
rect 5495 4503 5499 4559
rect 5499 4503 5555 4559
rect 5555 4503 5559 4559
rect 5495 4499 5559 4503
rect 5927 4559 5991 4563
rect 5927 4503 5931 4559
rect 5931 4503 5987 4559
rect 5987 4503 5991 4559
rect 5927 4499 5991 4503
rect 6271 4571 6335 4575
rect 6271 4515 6275 4571
rect 6275 4515 6331 4571
rect 6331 4515 6335 4571
rect 6271 4511 6335 4515
rect 6695 4571 6759 4575
rect 6695 4515 6699 4571
rect 6699 4515 6755 4571
rect 6755 4515 6759 4571
rect 6695 4511 6759 4515
rect 5023 4187 5087 4191
rect 5023 4131 5027 4187
rect 5027 4131 5083 4187
rect 5083 4131 5087 4187
rect 5023 4127 5087 4131
rect 5495 4187 5559 4191
rect 5495 4131 5499 4187
rect 5499 4131 5555 4187
rect 5555 4131 5559 4187
rect 5495 4127 5559 4131
rect 5927 4187 5991 4191
rect 5927 4131 5931 4187
rect 5931 4131 5987 4187
rect 5987 4131 5991 4187
rect 5927 4127 5991 4131
rect 6271 4175 6335 4179
rect 6271 4119 6275 4175
rect 6275 4119 6331 4175
rect 6331 4119 6335 4175
rect 6271 4115 6335 4119
rect 6695 4175 6759 4179
rect 6695 4119 6699 4175
rect 6699 4119 6755 4175
rect 6755 4119 6759 4175
rect 6695 4115 6759 4119
rect 5023 3769 5087 3773
rect 5023 3713 5027 3769
rect 5027 3713 5083 3769
rect 5083 3713 5087 3769
rect 5023 3709 5087 3713
rect 5495 3769 5559 3773
rect 5495 3713 5499 3769
rect 5499 3713 5555 3769
rect 5555 3713 5559 3769
rect 5495 3709 5559 3713
rect 5927 3769 5991 3773
rect 5927 3713 5931 3769
rect 5931 3713 5987 3769
rect 5987 3713 5991 3769
rect 5927 3709 5991 3713
rect 6271 3781 6335 3785
rect 6271 3725 6275 3781
rect 6275 3725 6331 3781
rect 6331 3725 6335 3781
rect 6271 3721 6335 3725
rect 6695 3781 6759 3785
rect 6695 3725 6699 3781
rect 6699 3725 6755 3781
rect 6755 3725 6759 3781
rect 6695 3721 6759 3725
rect 5023 3397 5087 3401
rect 5023 3341 5027 3397
rect 5027 3341 5083 3397
rect 5083 3341 5087 3397
rect 5023 3337 5087 3341
rect 5495 3397 5559 3401
rect 5495 3341 5499 3397
rect 5499 3341 5555 3397
rect 5555 3341 5559 3397
rect 5495 3337 5559 3341
rect 5927 3397 5991 3401
rect 5927 3341 5931 3397
rect 5931 3341 5987 3397
rect 5987 3341 5991 3397
rect 5927 3337 5991 3341
rect 6271 3385 6335 3389
rect 6271 3329 6275 3385
rect 6275 3329 6331 3385
rect 6331 3329 6335 3385
rect 6271 3325 6335 3329
rect 6695 3385 6759 3389
rect 6695 3329 6699 3385
rect 6699 3329 6755 3385
rect 6755 3329 6759 3385
rect 6695 3325 6759 3329
rect 5023 2979 5087 2983
rect 5023 2923 5027 2979
rect 5027 2923 5083 2979
rect 5083 2923 5087 2979
rect 5023 2919 5087 2923
rect 5495 2979 5559 2983
rect 5495 2923 5499 2979
rect 5499 2923 5555 2979
rect 5555 2923 5559 2979
rect 5495 2919 5559 2923
rect 5927 2979 5991 2983
rect 5927 2923 5931 2979
rect 5931 2923 5987 2979
rect 5987 2923 5991 2979
rect 5927 2919 5991 2923
rect 6271 2991 6335 2995
rect 6271 2935 6275 2991
rect 6275 2935 6331 2991
rect 6331 2935 6335 2991
rect 6271 2931 6335 2935
rect 6695 2991 6759 2995
rect 6695 2935 6699 2991
rect 6699 2935 6755 2991
rect 6755 2935 6759 2991
rect 6695 2931 6759 2935
rect 5023 2607 5087 2611
rect 5023 2551 5027 2607
rect 5027 2551 5083 2607
rect 5083 2551 5087 2607
rect 5023 2547 5087 2551
rect 5495 2607 5559 2611
rect 5495 2551 5499 2607
rect 5499 2551 5555 2607
rect 5555 2551 5559 2607
rect 5495 2547 5559 2551
rect 5927 2607 5991 2611
rect 5927 2551 5931 2607
rect 5931 2551 5987 2607
rect 5987 2551 5991 2607
rect 5927 2547 5991 2551
rect 6271 2595 6335 2599
rect 6271 2539 6275 2595
rect 6275 2539 6331 2595
rect 6331 2539 6335 2595
rect 6271 2535 6335 2539
rect 6695 2595 6759 2599
rect 6695 2539 6699 2595
rect 6699 2539 6755 2595
rect 6755 2539 6759 2595
rect 6695 2535 6759 2539
rect 5023 2189 5087 2193
rect 5023 2133 5027 2189
rect 5027 2133 5083 2189
rect 5083 2133 5087 2189
rect 5023 2129 5087 2133
rect 5495 2189 5559 2193
rect 5495 2133 5499 2189
rect 5499 2133 5555 2189
rect 5555 2133 5559 2189
rect 5495 2129 5559 2133
rect 5927 2189 5991 2193
rect 5927 2133 5931 2189
rect 5931 2133 5987 2189
rect 5987 2133 5991 2189
rect 5927 2129 5991 2133
rect 6271 2201 6335 2205
rect 6271 2145 6275 2201
rect 6275 2145 6331 2201
rect 6331 2145 6335 2201
rect 6271 2141 6335 2145
rect 6695 2201 6759 2205
rect 6695 2145 6699 2201
rect 6699 2145 6755 2201
rect 6755 2145 6759 2201
rect 6695 2141 6759 2145
rect 5023 1817 5087 1821
rect 5023 1761 5027 1817
rect 5027 1761 5083 1817
rect 5083 1761 5087 1817
rect 5023 1757 5087 1761
rect 5495 1817 5559 1821
rect 5495 1761 5499 1817
rect 5499 1761 5555 1817
rect 5555 1761 5559 1817
rect 5495 1757 5559 1761
rect 5927 1817 5991 1821
rect 5927 1761 5931 1817
rect 5931 1761 5987 1817
rect 5987 1761 5991 1817
rect 5927 1757 5991 1761
rect 6271 1805 6335 1809
rect 6271 1749 6275 1805
rect 6275 1749 6331 1805
rect 6331 1749 6335 1805
rect 6271 1745 6335 1749
rect 6695 1805 6759 1809
rect 6695 1749 6699 1805
rect 6699 1749 6755 1805
rect 6755 1749 6759 1805
rect 6695 1745 6759 1749
rect 5023 1399 5087 1403
rect 5023 1343 5027 1399
rect 5027 1343 5083 1399
rect 5083 1343 5087 1399
rect 5023 1339 5087 1343
rect 5495 1399 5559 1403
rect 5495 1343 5499 1399
rect 5499 1343 5555 1399
rect 5555 1343 5559 1399
rect 5495 1339 5559 1343
rect 5927 1399 5991 1403
rect 5927 1343 5931 1399
rect 5931 1343 5987 1399
rect 5987 1343 5991 1399
rect 5927 1339 5991 1343
rect 6271 1411 6335 1415
rect 6271 1355 6275 1411
rect 6275 1355 6331 1411
rect 6331 1355 6335 1411
rect 6271 1351 6335 1355
rect 6695 1411 6759 1415
rect 6695 1355 6699 1411
rect 6699 1355 6755 1411
rect 6755 1355 6759 1411
rect 6695 1351 6759 1355
rect 5023 1027 5087 1031
rect 5023 971 5027 1027
rect 5027 971 5083 1027
rect 5083 971 5087 1027
rect 5023 967 5087 971
rect 5495 1027 5559 1031
rect 5495 971 5499 1027
rect 5499 971 5555 1027
rect 5555 971 5559 1027
rect 5495 967 5559 971
rect 5927 1027 5991 1031
rect 5927 971 5931 1027
rect 5931 971 5987 1027
rect 5987 971 5991 1027
rect 5927 967 5991 971
rect 6271 1015 6335 1019
rect 6271 959 6275 1015
rect 6275 959 6331 1015
rect 6331 959 6335 1015
rect 6271 955 6335 959
rect 6695 1015 6759 1019
rect 6695 959 6699 1015
rect 6699 959 6755 1015
rect 6755 959 6759 1015
rect 6695 955 6759 959
rect 5023 609 5087 613
rect 5023 553 5027 609
rect 5027 553 5083 609
rect 5083 553 5087 609
rect 5023 549 5087 553
rect 5495 609 5559 613
rect 5495 553 5499 609
rect 5499 553 5555 609
rect 5555 553 5559 609
rect 5495 549 5559 553
rect 5927 609 5991 613
rect 5927 553 5931 609
rect 5931 553 5987 609
rect 5987 553 5991 609
rect 5927 549 5991 553
rect 6271 621 6335 625
rect 6271 565 6275 621
rect 6275 565 6331 621
rect 6331 565 6335 621
rect 6271 561 6335 565
rect 6695 621 6759 625
rect 6695 565 6699 621
rect 6699 565 6755 621
rect 6755 565 6759 621
rect 6695 561 6759 565
rect 5023 237 5087 241
rect 5023 181 5027 237
rect 5027 181 5083 237
rect 5083 181 5087 237
rect 5023 177 5087 181
rect 5495 237 5559 241
rect 5495 181 5499 237
rect 5499 181 5555 237
rect 5555 181 5559 237
rect 5495 177 5559 181
rect 5927 237 5991 241
rect 5927 181 5931 237
rect 5931 181 5987 237
rect 5987 181 5991 237
rect 5927 177 5991 181
rect 6271 225 6335 229
rect 6271 169 6275 225
rect 6275 169 6331 225
rect 6331 169 6335 225
rect 6271 165 6335 169
rect 6695 225 6759 229
rect 6695 169 6699 225
rect 6699 169 6755 225
rect 6755 169 6759 225
rect 6695 165 6759 169
<< metal4 >>
rect 5022 25103 5088 25341
rect 5022 25039 5023 25103
rect 5087 25039 5088 25103
rect 5022 24731 5088 25039
rect 5022 24667 5023 24731
rect 5087 24667 5088 24731
rect 5022 24313 5088 24667
rect 5022 24249 5023 24313
rect 5087 24249 5088 24313
rect 5022 23941 5088 24249
rect 5022 23877 5023 23941
rect 5087 23877 5088 23941
rect 5022 23523 5088 23877
rect 5022 23459 5023 23523
rect 5087 23459 5088 23523
rect 5022 23151 5088 23459
rect 5022 23087 5023 23151
rect 5087 23087 5088 23151
rect 5022 22733 5088 23087
rect 5022 22669 5023 22733
rect 5087 22669 5088 22733
rect 5022 22361 5088 22669
rect 5022 22297 5023 22361
rect 5087 22297 5088 22361
rect 5022 21943 5088 22297
rect 5022 21879 5023 21943
rect 5087 21879 5088 21943
rect 5022 21571 5088 21879
rect 5022 21507 5023 21571
rect 5087 21507 5088 21571
rect 5022 21153 5088 21507
rect 5022 21089 5023 21153
rect 5087 21089 5088 21153
rect 5022 20781 5088 21089
rect 5022 20717 5023 20781
rect 5087 20717 5088 20781
rect 5022 20363 5088 20717
rect 5022 20299 5023 20363
rect 5087 20299 5088 20363
rect 5022 19991 5088 20299
rect 5022 19927 5023 19991
rect 5087 19927 5088 19991
rect 5022 19573 5088 19927
rect 5022 19509 5023 19573
rect 5087 19509 5088 19573
rect 5022 19201 5088 19509
rect 5022 19137 5023 19201
rect 5087 19137 5088 19201
rect 5022 18783 5088 19137
rect 5022 18719 5023 18783
rect 5087 18719 5088 18783
rect 5022 18411 5088 18719
rect 5022 18347 5023 18411
rect 5087 18347 5088 18411
rect 5022 17993 5088 18347
rect 5022 17929 5023 17993
rect 5087 17929 5088 17993
rect 5022 17621 5088 17929
rect 5022 17557 5023 17621
rect 5087 17557 5088 17621
rect 5022 17203 5088 17557
rect 5022 17139 5023 17203
rect 5087 17139 5088 17203
rect 5022 16831 5088 17139
rect 5022 16767 5023 16831
rect 5087 16767 5088 16831
rect 5022 16413 5088 16767
rect 5022 16349 5023 16413
rect 5087 16349 5088 16413
rect 5022 16041 5088 16349
rect 5022 15977 5023 16041
rect 5087 15977 5088 16041
rect 5022 15623 5088 15977
rect 5022 15559 5023 15623
rect 5087 15559 5088 15623
rect 5022 15251 5088 15559
rect 5022 15187 5023 15251
rect 5087 15187 5088 15251
rect 5022 14833 5088 15187
rect 5022 14769 5023 14833
rect 5087 14769 5088 14833
rect 5022 14461 5088 14769
rect 5022 14397 5023 14461
rect 5087 14397 5088 14461
rect 5022 14043 5088 14397
rect 5022 13979 5023 14043
rect 5087 13979 5088 14043
rect 5022 13671 5088 13979
rect 5022 13607 5023 13671
rect 5087 13607 5088 13671
rect 5022 13253 5088 13607
rect 5022 13189 5023 13253
rect 5087 13189 5088 13253
rect 5022 12881 5088 13189
rect 5022 12817 5023 12881
rect 5087 12817 5088 12881
rect 5022 12463 5088 12817
rect 5022 12399 5023 12463
rect 5087 12399 5088 12463
rect 5022 12091 5088 12399
rect 5022 12027 5023 12091
rect 5087 12027 5088 12091
rect 5022 11673 5088 12027
rect 5022 11609 5023 11673
rect 5087 11609 5088 11673
rect 5022 11301 5088 11609
rect 5022 11237 5023 11301
rect 5087 11237 5088 11301
rect 5022 10883 5088 11237
rect 5022 10819 5023 10883
rect 5087 10819 5088 10883
rect 5022 10511 5088 10819
rect 5022 10447 5023 10511
rect 5087 10447 5088 10511
rect 5022 10093 5088 10447
rect 5022 10029 5023 10093
rect 5087 10029 5088 10093
rect 5022 9721 5088 10029
rect 5022 9657 5023 9721
rect 5087 9657 5088 9721
rect 5022 9303 5088 9657
rect 5022 9239 5023 9303
rect 5087 9239 5088 9303
rect 5022 8931 5088 9239
rect 5022 8867 5023 8931
rect 5087 8867 5088 8931
rect 5022 8513 5088 8867
rect 5022 8449 5023 8513
rect 5087 8449 5088 8513
rect 5022 8141 5088 8449
rect 5022 8077 5023 8141
rect 5087 8077 5088 8141
rect 5022 7723 5088 8077
rect 5022 7659 5023 7723
rect 5087 7659 5088 7723
rect 5022 7351 5088 7659
rect 5022 7287 5023 7351
rect 5087 7287 5088 7351
rect 5022 6933 5088 7287
rect 5022 6869 5023 6933
rect 5087 6869 5088 6933
rect 5022 6561 5088 6869
rect 5022 6497 5023 6561
rect 5087 6497 5088 6561
rect 5022 6143 5088 6497
rect 5022 6079 5023 6143
rect 5087 6079 5088 6143
rect 5022 5771 5088 6079
rect 5022 5707 5023 5771
rect 5087 5707 5088 5771
rect 5022 5353 5088 5707
rect 5022 5289 5023 5353
rect 5087 5289 5088 5353
rect 5022 4981 5088 5289
rect 5022 4917 5023 4981
rect 5087 4917 5088 4981
rect 5022 4563 5088 4917
rect 5022 4499 5023 4563
rect 5087 4499 5088 4563
rect 5022 4191 5088 4499
rect 5022 4127 5023 4191
rect 5087 4127 5088 4191
rect 5022 3773 5088 4127
rect 5022 3709 5023 3773
rect 5087 3709 5088 3773
rect 5022 3401 5088 3709
rect 5022 3337 5023 3401
rect 5087 3337 5088 3401
rect 5022 2983 5088 3337
rect 5022 2919 5023 2983
rect 5087 2919 5088 2983
rect 5022 2611 5088 2919
rect 5022 2547 5023 2611
rect 5087 2547 5088 2611
rect 5022 2193 5088 2547
rect 5022 2129 5023 2193
rect 5087 2129 5088 2193
rect 5022 1821 5088 2129
rect 5022 1757 5023 1821
rect 5087 1757 5088 1821
rect 5022 1403 5088 1757
rect 5022 1339 5023 1403
rect 5087 1339 5088 1403
rect 5022 1031 5088 1339
rect 5022 967 5023 1031
rect 5087 967 5088 1031
rect 5022 613 5088 967
rect 5022 549 5023 613
rect 5087 549 5088 613
rect 5022 241 5088 549
rect 5022 177 5023 241
rect 5087 177 5088 241
rect 5022 -33 5088 177
rect 5494 25103 5560 25341
rect 5494 25039 5495 25103
rect 5559 25039 5560 25103
rect 5494 24731 5560 25039
rect 5494 24667 5495 24731
rect 5559 24667 5560 24731
rect 5494 24313 5560 24667
rect 5494 24249 5495 24313
rect 5559 24249 5560 24313
rect 5494 23941 5560 24249
rect 5494 23877 5495 23941
rect 5559 23877 5560 23941
rect 5494 23523 5560 23877
rect 5494 23459 5495 23523
rect 5559 23459 5560 23523
rect 5494 23151 5560 23459
rect 5494 23087 5495 23151
rect 5559 23087 5560 23151
rect 5494 22733 5560 23087
rect 5494 22669 5495 22733
rect 5559 22669 5560 22733
rect 5494 22361 5560 22669
rect 5494 22297 5495 22361
rect 5559 22297 5560 22361
rect 5494 21943 5560 22297
rect 5494 21879 5495 21943
rect 5559 21879 5560 21943
rect 5494 21571 5560 21879
rect 5494 21507 5495 21571
rect 5559 21507 5560 21571
rect 5494 21153 5560 21507
rect 5494 21089 5495 21153
rect 5559 21089 5560 21153
rect 5494 20781 5560 21089
rect 5494 20717 5495 20781
rect 5559 20717 5560 20781
rect 5494 20363 5560 20717
rect 5494 20299 5495 20363
rect 5559 20299 5560 20363
rect 5494 19991 5560 20299
rect 5494 19927 5495 19991
rect 5559 19927 5560 19991
rect 5494 19573 5560 19927
rect 5494 19509 5495 19573
rect 5559 19509 5560 19573
rect 5494 19201 5560 19509
rect 5494 19137 5495 19201
rect 5559 19137 5560 19201
rect 5494 18783 5560 19137
rect 5494 18719 5495 18783
rect 5559 18719 5560 18783
rect 5494 18411 5560 18719
rect 5494 18347 5495 18411
rect 5559 18347 5560 18411
rect 5494 17993 5560 18347
rect 5494 17929 5495 17993
rect 5559 17929 5560 17993
rect 5494 17621 5560 17929
rect 5494 17557 5495 17621
rect 5559 17557 5560 17621
rect 5494 17203 5560 17557
rect 5494 17139 5495 17203
rect 5559 17139 5560 17203
rect 5494 16831 5560 17139
rect 5494 16767 5495 16831
rect 5559 16767 5560 16831
rect 5494 16413 5560 16767
rect 5494 16349 5495 16413
rect 5559 16349 5560 16413
rect 5494 16041 5560 16349
rect 5494 15977 5495 16041
rect 5559 15977 5560 16041
rect 5494 15623 5560 15977
rect 5494 15559 5495 15623
rect 5559 15559 5560 15623
rect 5494 15251 5560 15559
rect 5494 15187 5495 15251
rect 5559 15187 5560 15251
rect 5494 14833 5560 15187
rect 5494 14769 5495 14833
rect 5559 14769 5560 14833
rect 5494 14461 5560 14769
rect 5494 14397 5495 14461
rect 5559 14397 5560 14461
rect 5494 14043 5560 14397
rect 5494 13979 5495 14043
rect 5559 13979 5560 14043
rect 5494 13671 5560 13979
rect 5494 13607 5495 13671
rect 5559 13607 5560 13671
rect 5494 13253 5560 13607
rect 5494 13189 5495 13253
rect 5559 13189 5560 13253
rect 5494 12881 5560 13189
rect 5494 12817 5495 12881
rect 5559 12817 5560 12881
rect 5494 12463 5560 12817
rect 5494 12399 5495 12463
rect 5559 12399 5560 12463
rect 5494 12091 5560 12399
rect 5494 12027 5495 12091
rect 5559 12027 5560 12091
rect 5494 11673 5560 12027
rect 5494 11609 5495 11673
rect 5559 11609 5560 11673
rect 5494 11301 5560 11609
rect 5494 11237 5495 11301
rect 5559 11237 5560 11301
rect 5494 10883 5560 11237
rect 5494 10819 5495 10883
rect 5559 10819 5560 10883
rect 5494 10511 5560 10819
rect 5494 10447 5495 10511
rect 5559 10447 5560 10511
rect 5494 10093 5560 10447
rect 5494 10029 5495 10093
rect 5559 10029 5560 10093
rect 5494 9721 5560 10029
rect 5494 9657 5495 9721
rect 5559 9657 5560 9721
rect 5494 9303 5560 9657
rect 5494 9239 5495 9303
rect 5559 9239 5560 9303
rect 5494 8931 5560 9239
rect 5494 8867 5495 8931
rect 5559 8867 5560 8931
rect 5494 8513 5560 8867
rect 5494 8449 5495 8513
rect 5559 8449 5560 8513
rect 5494 8141 5560 8449
rect 5494 8077 5495 8141
rect 5559 8077 5560 8141
rect 5494 7723 5560 8077
rect 5494 7659 5495 7723
rect 5559 7659 5560 7723
rect 5494 7351 5560 7659
rect 5494 7287 5495 7351
rect 5559 7287 5560 7351
rect 5494 6933 5560 7287
rect 5494 6869 5495 6933
rect 5559 6869 5560 6933
rect 5494 6561 5560 6869
rect 5494 6497 5495 6561
rect 5559 6497 5560 6561
rect 5494 6143 5560 6497
rect 5494 6079 5495 6143
rect 5559 6079 5560 6143
rect 5494 5771 5560 6079
rect 5494 5707 5495 5771
rect 5559 5707 5560 5771
rect 5494 5353 5560 5707
rect 5494 5289 5495 5353
rect 5559 5289 5560 5353
rect 5494 4981 5560 5289
rect 5494 4917 5495 4981
rect 5559 4917 5560 4981
rect 5494 4563 5560 4917
rect 5494 4499 5495 4563
rect 5559 4499 5560 4563
rect 5494 4191 5560 4499
rect 5494 4127 5495 4191
rect 5559 4127 5560 4191
rect 5494 3773 5560 4127
rect 5494 3709 5495 3773
rect 5559 3709 5560 3773
rect 5494 3401 5560 3709
rect 5494 3337 5495 3401
rect 5559 3337 5560 3401
rect 5494 2983 5560 3337
rect 5494 2919 5495 2983
rect 5559 2919 5560 2983
rect 5494 2611 5560 2919
rect 5494 2547 5495 2611
rect 5559 2547 5560 2611
rect 5494 2193 5560 2547
rect 5494 2129 5495 2193
rect 5559 2129 5560 2193
rect 5494 1821 5560 2129
rect 5494 1757 5495 1821
rect 5559 1757 5560 1821
rect 5494 1403 5560 1757
rect 5494 1339 5495 1403
rect 5559 1339 5560 1403
rect 5494 1031 5560 1339
rect 5494 967 5495 1031
rect 5559 967 5560 1031
rect 5494 613 5560 967
rect 5494 549 5495 613
rect 5559 549 5560 613
rect 5494 241 5560 549
rect 5494 177 5495 241
rect 5559 177 5560 241
rect 5494 -33 5560 177
rect 5926 25103 5992 25341
rect 5926 25039 5927 25103
rect 5991 25039 5992 25103
rect 5926 24731 5992 25039
rect 5926 24667 5927 24731
rect 5991 24667 5992 24731
rect 5926 24313 5992 24667
rect 5926 24249 5927 24313
rect 5991 24249 5992 24313
rect 5926 23941 5992 24249
rect 5926 23877 5927 23941
rect 5991 23877 5992 23941
rect 5926 23523 5992 23877
rect 5926 23459 5927 23523
rect 5991 23459 5992 23523
rect 5926 23151 5992 23459
rect 5926 23087 5927 23151
rect 5991 23087 5992 23151
rect 5926 22733 5992 23087
rect 5926 22669 5927 22733
rect 5991 22669 5992 22733
rect 5926 22361 5992 22669
rect 5926 22297 5927 22361
rect 5991 22297 5992 22361
rect 5926 21943 5992 22297
rect 5926 21879 5927 21943
rect 5991 21879 5992 21943
rect 5926 21571 5992 21879
rect 5926 21507 5927 21571
rect 5991 21507 5992 21571
rect 5926 21153 5992 21507
rect 5926 21089 5927 21153
rect 5991 21089 5992 21153
rect 5926 20781 5992 21089
rect 5926 20717 5927 20781
rect 5991 20717 5992 20781
rect 5926 20363 5992 20717
rect 5926 20299 5927 20363
rect 5991 20299 5992 20363
rect 5926 19991 5992 20299
rect 5926 19927 5927 19991
rect 5991 19927 5992 19991
rect 5926 19573 5992 19927
rect 5926 19509 5927 19573
rect 5991 19509 5992 19573
rect 5926 19201 5992 19509
rect 5926 19137 5927 19201
rect 5991 19137 5992 19201
rect 5926 18783 5992 19137
rect 5926 18719 5927 18783
rect 5991 18719 5992 18783
rect 5926 18411 5992 18719
rect 5926 18347 5927 18411
rect 5991 18347 5992 18411
rect 5926 17993 5992 18347
rect 5926 17929 5927 17993
rect 5991 17929 5992 17993
rect 5926 17621 5992 17929
rect 5926 17557 5927 17621
rect 5991 17557 5992 17621
rect 5926 17203 5992 17557
rect 5926 17139 5927 17203
rect 5991 17139 5992 17203
rect 5926 16831 5992 17139
rect 5926 16767 5927 16831
rect 5991 16767 5992 16831
rect 5926 16413 5992 16767
rect 5926 16349 5927 16413
rect 5991 16349 5992 16413
rect 5926 16041 5992 16349
rect 5926 15977 5927 16041
rect 5991 15977 5992 16041
rect 5926 15623 5992 15977
rect 5926 15559 5927 15623
rect 5991 15559 5992 15623
rect 5926 15251 5992 15559
rect 5926 15187 5927 15251
rect 5991 15187 5992 15251
rect 5926 14833 5992 15187
rect 5926 14769 5927 14833
rect 5991 14769 5992 14833
rect 5926 14461 5992 14769
rect 5926 14397 5927 14461
rect 5991 14397 5992 14461
rect 5926 14043 5992 14397
rect 5926 13979 5927 14043
rect 5991 13979 5992 14043
rect 5926 13671 5992 13979
rect 5926 13607 5927 13671
rect 5991 13607 5992 13671
rect 5926 13253 5992 13607
rect 5926 13189 5927 13253
rect 5991 13189 5992 13253
rect 5926 12881 5992 13189
rect 5926 12817 5927 12881
rect 5991 12817 5992 12881
rect 5926 12463 5992 12817
rect 5926 12399 5927 12463
rect 5991 12399 5992 12463
rect 5926 12091 5992 12399
rect 5926 12027 5927 12091
rect 5991 12027 5992 12091
rect 5926 11673 5992 12027
rect 5926 11609 5927 11673
rect 5991 11609 5992 11673
rect 5926 11301 5992 11609
rect 5926 11237 5927 11301
rect 5991 11237 5992 11301
rect 5926 10883 5992 11237
rect 5926 10819 5927 10883
rect 5991 10819 5992 10883
rect 5926 10511 5992 10819
rect 5926 10447 5927 10511
rect 5991 10447 5992 10511
rect 5926 10093 5992 10447
rect 5926 10029 5927 10093
rect 5991 10029 5992 10093
rect 5926 9721 5992 10029
rect 5926 9657 5927 9721
rect 5991 9657 5992 9721
rect 5926 9303 5992 9657
rect 5926 9239 5927 9303
rect 5991 9239 5992 9303
rect 5926 8931 5992 9239
rect 5926 8867 5927 8931
rect 5991 8867 5992 8931
rect 5926 8513 5992 8867
rect 5926 8449 5927 8513
rect 5991 8449 5992 8513
rect 5926 8141 5992 8449
rect 5926 8077 5927 8141
rect 5991 8077 5992 8141
rect 5926 7723 5992 8077
rect 5926 7659 5927 7723
rect 5991 7659 5992 7723
rect 5926 7351 5992 7659
rect 5926 7287 5927 7351
rect 5991 7287 5992 7351
rect 5926 6933 5992 7287
rect 5926 6869 5927 6933
rect 5991 6869 5992 6933
rect 5926 6561 5992 6869
rect 5926 6497 5927 6561
rect 5991 6497 5992 6561
rect 5926 6143 5992 6497
rect 5926 6079 5927 6143
rect 5991 6079 5992 6143
rect 5926 5771 5992 6079
rect 5926 5707 5927 5771
rect 5991 5707 5992 5771
rect 5926 5353 5992 5707
rect 5926 5289 5927 5353
rect 5991 5289 5992 5353
rect 5926 4981 5992 5289
rect 5926 4917 5927 4981
rect 5991 4917 5992 4981
rect 5926 4563 5992 4917
rect 5926 4499 5927 4563
rect 5991 4499 5992 4563
rect 5926 4191 5992 4499
rect 5926 4127 5927 4191
rect 5991 4127 5992 4191
rect 5926 3773 5992 4127
rect 5926 3709 5927 3773
rect 5991 3709 5992 3773
rect 5926 3401 5992 3709
rect 5926 3337 5927 3401
rect 5991 3337 5992 3401
rect 5926 2983 5992 3337
rect 5926 2919 5927 2983
rect 5991 2919 5992 2983
rect 5926 2611 5992 2919
rect 5926 2547 5927 2611
rect 5991 2547 5992 2611
rect 5926 2193 5992 2547
rect 5926 2129 5927 2193
rect 5991 2129 5992 2193
rect 5926 1821 5992 2129
rect 5926 1757 5927 1821
rect 5991 1757 5992 1821
rect 5926 1403 5992 1757
rect 5926 1339 5927 1403
rect 5991 1339 5992 1403
rect 5926 1031 5992 1339
rect 5926 967 5927 1031
rect 5991 967 5992 1031
rect 5926 613 5992 967
rect 5926 549 5927 613
rect 5991 549 5992 613
rect 5926 241 5992 549
rect 5926 177 5927 241
rect 5991 177 5992 241
rect 5926 -33 5992 177
rect 6270 25115 6336 25341
rect 6270 25051 6271 25115
rect 6335 25051 6336 25115
rect 6270 24719 6336 25051
rect 6270 24655 6271 24719
rect 6335 24655 6336 24719
rect 6270 24325 6336 24655
rect 6270 24261 6271 24325
rect 6335 24261 6336 24325
rect 6270 23929 6336 24261
rect 6270 23865 6271 23929
rect 6335 23865 6336 23929
rect 6270 23535 6336 23865
rect 6270 23471 6271 23535
rect 6335 23471 6336 23535
rect 6270 23139 6336 23471
rect 6270 23075 6271 23139
rect 6335 23075 6336 23139
rect 6270 22745 6336 23075
rect 6270 22681 6271 22745
rect 6335 22681 6336 22745
rect 6270 22349 6336 22681
rect 6270 22285 6271 22349
rect 6335 22285 6336 22349
rect 6270 21955 6336 22285
rect 6270 21891 6271 21955
rect 6335 21891 6336 21955
rect 6270 21559 6336 21891
rect 6270 21495 6271 21559
rect 6335 21495 6336 21559
rect 6270 21165 6336 21495
rect 6270 21101 6271 21165
rect 6335 21101 6336 21165
rect 6270 20769 6336 21101
rect 6270 20705 6271 20769
rect 6335 20705 6336 20769
rect 6270 20375 6336 20705
rect 6270 20311 6271 20375
rect 6335 20311 6336 20375
rect 6270 19979 6336 20311
rect 6270 19915 6271 19979
rect 6335 19915 6336 19979
rect 6270 19585 6336 19915
rect 6270 19521 6271 19585
rect 6335 19521 6336 19585
rect 6270 19189 6336 19521
rect 6270 19125 6271 19189
rect 6335 19125 6336 19189
rect 6270 18795 6336 19125
rect 6270 18731 6271 18795
rect 6335 18731 6336 18795
rect 6270 18399 6336 18731
rect 6270 18335 6271 18399
rect 6335 18335 6336 18399
rect 6270 18005 6336 18335
rect 6270 17941 6271 18005
rect 6335 17941 6336 18005
rect 6270 17609 6336 17941
rect 6270 17545 6271 17609
rect 6335 17545 6336 17609
rect 6270 17215 6336 17545
rect 6270 17151 6271 17215
rect 6335 17151 6336 17215
rect 6270 16819 6336 17151
rect 6270 16755 6271 16819
rect 6335 16755 6336 16819
rect 6270 16425 6336 16755
rect 6270 16361 6271 16425
rect 6335 16361 6336 16425
rect 6270 16029 6336 16361
rect 6270 15965 6271 16029
rect 6335 15965 6336 16029
rect 6270 15635 6336 15965
rect 6270 15571 6271 15635
rect 6335 15571 6336 15635
rect 6270 15239 6336 15571
rect 6270 15175 6271 15239
rect 6335 15175 6336 15239
rect 6270 14845 6336 15175
rect 6270 14781 6271 14845
rect 6335 14781 6336 14845
rect 6270 14449 6336 14781
rect 6270 14385 6271 14449
rect 6335 14385 6336 14449
rect 6270 14055 6336 14385
rect 6270 13991 6271 14055
rect 6335 13991 6336 14055
rect 6270 13659 6336 13991
rect 6270 13595 6271 13659
rect 6335 13595 6336 13659
rect 6270 13265 6336 13595
rect 6270 13201 6271 13265
rect 6335 13201 6336 13265
rect 6270 12869 6336 13201
rect 6270 12805 6271 12869
rect 6335 12805 6336 12869
rect 6270 12475 6336 12805
rect 6270 12411 6271 12475
rect 6335 12411 6336 12475
rect 6270 12079 6336 12411
rect 6270 12015 6271 12079
rect 6335 12015 6336 12079
rect 6270 11685 6336 12015
rect 6270 11621 6271 11685
rect 6335 11621 6336 11685
rect 6270 11289 6336 11621
rect 6270 11225 6271 11289
rect 6335 11225 6336 11289
rect 6270 10895 6336 11225
rect 6270 10831 6271 10895
rect 6335 10831 6336 10895
rect 6270 10499 6336 10831
rect 6270 10435 6271 10499
rect 6335 10435 6336 10499
rect 6270 10105 6336 10435
rect 6270 10041 6271 10105
rect 6335 10041 6336 10105
rect 6270 9709 6336 10041
rect 6270 9645 6271 9709
rect 6335 9645 6336 9709
rect 6270 9315 6336 9645
rect 6270 9251 6271 9315
rect 6335 9251 6336 9315
rect 6270 8919 6336 9251
rect 6270 8855 6271 8919
rect 6335 8855 6336 8919
rect 6270 8525 6336 8855
rect 6270 8461 6271 8525
rect 6335 8461 6336 8525
rect 6270 8129 6336 8461
rect 6270 8065 6271 8129
rect 6335 8065 6336 8129
rect 6270 7735 6336 8065
rect 6270 7671 6271 7735
rect 6335 7671 6336 7735
rect 6270 7339 6336 7671
rect 6270 7275 6271 7339
rect 6335 7275 6336 7339
rect 6270 6945 6336 7275
rect 6270 6881 6271 6945
rect 6335 6881 6336 6945
rect 6270 6549 6336 6881
rect 6270 6485 6271 6549
rect 6335 6485 6336 6549
rect 6270 6155 6336 6485
rect 6270 6091 6271 6155
rect 6335 6091 6336 6155
rect 6270 5759 6336 6091
rect 6270 5695 6271 5759
rect 6335 5695 6336 5759
rect 6270 5365 6336 5695
rect 6270 5301 6271 5365
rect 6335 5301 6336 5365
rect 6270 4969 6336 5301
rect 6270 4905 6271 4969
rect 6335 4905 6336 4969
rect 6270 4575 6336 4905
rect 6270 4511 6271 4575
rect 6335 4511 6336 4575
rect 6270 4179 6336 4511
rect 6270 4115 6271 4179
rect 6335 4115 6336 4179
rect 6270 3785 6336 4115
rect 6270 3721 6271 3785
rect 6335 3721 6336 3785
rect 6270 3389 6336 3721
rect 6270 3325 6271 3389
rect 6335 3325 6336 3389
rect 6270 2995 6336 3325
rect 6270 2931 6271 2995
rect 6335 2931 6336 2995
rect 6270 2599 6336 2931
rect 6270 2535 6271 2599
rect 6335 2535 6336 2599
rect 6270 2205 6336 2535
rect 6270 2141 6271 2205
rect 6335 2141 6336 2205
rect 6270 1809 6336 2141
rect 6270 1745 6271 1809
rect 6335 1745 6336 1809
rect 6270 1415 6336 1745
rect 6270 1351 6271 1415
rect 6335 1351 6336 1415
rect 6270 1019 6336 1351
rect 6270 955 6271 1019
rect 6335 955 6336 1019
rect 6270 625 6336 955
rect 6270 561 6271 625
rect 6335 561 6336 625
rect 6270 229 6336 561
rect 6270 165 6271 229
rect 6335 165 6336 229
rect 6270 -33 6336 165
rect 6694 25115 6760 25341
rect 6694 25051 6695 25115
rect 6759 25051 6760 25115
rect 6694 24719 6760 25051
rect 6694 24655 6695 24719
rect 6759 24655 6760 24719
rect 6694 24325 6760 24655
rect 6694 24261 6695 24325
rect 6759 24261 6760 24325
rect 6694 23929 6760 24261
rect 6694 23865 6695 23929
rect 6759 23865 6760 23929
rect 6694 23535 6760 23865
rect 6694 23471 6695 23535
rect 6759 23471 6760 23535
rect 6694 23139 6760 23471
rect 6694 23075 6695 23139
rect 6759 23075 6760 23139
rect 6694 22745 6760 23075
rect 6694 22681 6695 22745
rect 6759 22681 6760 22745
rect 6694 22349 6760 22681
rect 6694 22285 6695 22349
rect 6759 22285 6760 22349
rect 6694 21955 6760 22285
rect 6694 21891 6695 21955
rect 6759 21891 6760 21955
rect 6694 21559 6760 21891
rect 6694 21495 6695 21559
rect 6759 21495 6760 21559
rect 6694 21165 6760 21495
rect 6694 21101 6695 21165
rect 6759 21101 6760 21165
rect 6694 20769 6760 21101
rect 6694 20705 6695 20769
rect 6759 20705 6760 20769
rect 6694 20375 6760 20705
rect 6694 20311 6695 20375
rect 6759 20311 6760 20375
rect 6694 19979 6760 20311
rect 6694 19915 6695 19979
rect 6759 19915 6760 19979
rect 6694 19585 6760 19915
rect 6694 19521 6695 19585
rect 6759 19521 6760 19585
rect 6694 19189 6760 19521
rect 6694 19125 6695 19189
rect 6759 19125 6760 19189
rect 6694 18795 6760 19125
rect 6694 18731 6695 18795
rect 6759 18731 6760 18795
rect 6694 18399 6760 18731
rect 6694 18335 6695 18399
rect 6759 18335 6760 18399
rect 6694 18005 6760 18335
rect 6694 17941 6695 18005
rect 6759 17941 6760 18005
rect 6694 17609 6760 17941
rect 6694 17545 6695 17609
rect 6759 17545 6760 17609
rect 6694 17215 6760 17545
rect 6694 17151 6695 17215
rect 6759 17151 6760 17215
rect 6694 16819 6760 17151
rect 6694 16755 6695 16819
rect 6759 16755 6760 16819
rect 6694 16425 6760 16755
rect 6694 16361 6695 16425
rect 6759 16361 6760 16425
rect 6694 16029 6760 16361
rect 6694 15965 6695 16029
rect 6759 15965 6760 16029
rect 6694 15635 6760 15965
rect 6694 15571 6695 15635
rect 6759 15571 6760 15635
rect 6694 15239 6760 15571
rect 6694 15175 6695 15239
rect 6759 15175 6760 15239
rect 6694 14845 6760 15175
rect 6694 14781 6695 14845
rect 6759 14781 6760 14845
rect 6694 14449 6760 14781
rect 6694 14385 6695 14449
rect 6759 14385 6760 14449
rect 6694 14055 6760 14385
rect 6694 13991 6695 14055
rect 6759 13991 6760 14055
rect 6694 13659 6760 13991
rect 6694 13595 6695 13659
rect 6759 13595 6760 13659
rect 6694 13265 6760 13595
rect 6694 13201 6695 13265
rect 6759 13201 6760 13265
rect 6694 12869 6760 13201
rect 6694 12805 6695 12869
rect 6759 12805 6760 12869
rect 6694 12475 6760 12805
rect 6694 12411 6695 12475
rect 6759 12411 6760 12475
rect 6694 12079 6760 12411
rect 6694 12015 6695 12079
rect 6759 12015 6760 12079
rect 6694 11685 6760 12015
rect 6694 11621 6695 11685
rect 6759 11621 6760 11685
rect 6694 11289 6760 11621
rect 6694 11225 6695 11289
rect 6759 11225 6760 11289
rect 6694 10895 6760 11225
rect 6694 10831 6695 10895
rect 6759 10831 6760 10895
rect 6694 10499 6760 10831
rect 6694 10435 6695 10499
rect 6759 10435 6760 10499
rect 6694 10105 6760 10435
rect 6694 10041 6695 10105
rect 6759 10041 6760 10105
rect 6694 9709 6760 10041
rect 6694 9645 6695 9709
rect 6759 9645 6760 9709
rect 6694 9315 6760 9645
rect 6694 9251 6695 9315
rect 6759 9251 6760 9315
rect 6694 8919 6760 9251
rect 6694 8855 6695 8919
rect 6759 8855 6760 8919
rect 6694 8525 6760 8855
rect 6694 8461 6695 8525
rect 6759 8461 6760 8525
rect 6694 8129 6760 8461
rect 6694 8065 6695 8129
rect 6759 8065 6760 8129
rect 6694 7735 6760 8065
rect 6694 7671 6695 7735
rect 6759 7671 6760 7735
rect 6694 7339 6760 7671
rect 6694 7275 6695 7339
rect 6759 7275 6760 7339
rect 6694 6945 6760 7275
rect 6694 6881 6695 6945
rect 6759 6881 6760 6945
rect 6694 6549 6760 6881
rect 6694 6485 6695 6549
rect 6759 6485 6760 6549
rect 6694 6155 6760 6485
rect 6694 6091 6695 6155
rect 6759 6091 6760 6155
rect 6694 5759 6760 6091
rect 6694 5695 6695 5759
rect 6759 5695 6760 5759
rect 6694 5365 6760 5695
rect 6694 5301 6695 5365
rect 6759 5301 6760 5365
rect 6694 4969 6760 5301
rect 6694 4905 6695 4969
rect 6759 4905 6760 4969
rect 6694 4575 6760 4905
rect 6694 4511 6695 4575
rect 6759 4511 6760 4575
rect 6694 4179 6760 4511
rect 6694 4115 6695 4179
rect 6759 4115 6760 4179
rect 6694 3785 6760 4115
rect 6694 3721 6695 3785
rect 6759 3721 6760 3785
rect 6694 3389 6760 3721
rect 6694 3325 6695 3389
rect 6759 3325 6760 3389
rect 6694 2995 6760 3325
rect 6694 2931 6695 2995
rect 6759 2931 6760 2995
rect 6694 2599 6760 2931
rect 6694 2535 6695 2599
rect 6759 2535 6760 2599
rect 6694 2205 6760 2535
rect 6694 2141 6695 2205
rect 6759 2141 6760 2205
rect 6694 1809 6760 2141
rect 6694 1745 6695 1809
rect 6759 1745 6760 1809
rect 6694 1415 6760 1745
rect 6694 1351 6695 1415
rect 6759 1351 6760 1415
rect 6694 1019 6760 1351
rect 6694 955 6695 1019
rect 6759 955 6760 1019
rect 6694 625 6760 955
rect 6694 561 6695 625
rect 6759 561 6760 625
rect 6694 229 6760 561
rect 6694 165 6695 229
rect 6759 165 6760 229
rect 6694 -33 6760 165
use subbyte2_and3_dec  subbyte2_and3_dec_0
timestamp 1543373569
transform 1 0 4807 0 -1 25280
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_1
timestamp 1543373569
transform 1 0 4807 0 1 24490
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_2
timestamp 1543373569
transform 1 0 4807 0 -1 24490
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_3
timestamp 1543373569
transform 1 0 4807 0 1 23700
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_4
timestamp 1543373569
transform 1 0 4807 0 -1 23700
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_5
timestamp 1543373569
transform 1 0 4807 0 1 22910
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_6
timestamp 1543373569
transform 1 0 4807 0 -1 22910
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_7
timestamp 1543373569
transform 1 0 4807 0 1 22120
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_8
timestamp 1543373569
transform 1 0 4807 0 -1 22120
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_9
timestamp 1543373569
transform 1 0 4807 0 1 21330
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_10
timestamp 1543373569
transform 1 0 4807 0 -1 21330
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_11
timestamp 1543373569
transform 1 0 4807 0 1 20540
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_12
timestamp 1543373569
transform 1 0 4807 0 -1 20540
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_13
timestamp 1543373569
transform 1 0 4807 0 1 19750
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_14
timestamp 1543373569
transform 1 0 4807 0 -1 19750
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_15
timestamp 1543373569
transform 1 0 4807 0 1 18960
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_16
timestamp 1543373569
transform 1 0 4807 0 -1 18960
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_17
timestamp 1543373569
transform 1 0 4807 0 1 18170
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_18
timestamp 1543373569
transform 1 0 4807 0 -1 18170
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_19
timestamp 1543373569
transform 1 0 4807 0 1 17380
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_20
timestamp 1543373569
transform 1 0 4807 0 -1 17380
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_21
timestamp 1543373569
transform 1 0 4807 0 1 16590
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_22
timestamp 1543373569
transform 1 0 4807 0 -1 16590
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_23
timestamp 1543373569
transform 1 0 4807 0 1 15800
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_24
timestamp 1543373569
transform 1 0 4807 0 -1 15800
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_25
timestamp 1543373569
transform 1 0 4807 0 1 15010
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_26
timestamp 1543373569
transform 1 0 4807 0 -1 15010
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_27
timestamp 1543373569
transform 1 0 4807 0 1 14220
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_28
timestamp 1543373569
transform 1 0 4807 0 -1 14220
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_29
timestamp 1543373569
transform 1 0 4807 0 1 13430
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_30
timestamp 1543373569
transform 1 0 4807 0 -1 13430
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_31
timestamp 1543373569
transform 1 0 4807 0 1 12640
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_32
timestamp 1543373569
transform 1 0 4807 0 -1 12640
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_33
timestamp 1543373569
transform 1 0 4807 0 1 11850
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_34
timestamp 1543373569
transform 1 0 4807 0 -1 11850
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_35
timestamp 1543373569
transform 1 0 4807 0 1 11060
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_36
timestamp 1543373569
transform 1 0 4807 0 -1 11060
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_37
timestamp 1543373569
transform 1 0 4807 0 1 10270
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_38
timestamp 1543373569
transform 1 0 4807 0 -1 10270
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_39
timestamp 1543373569
transform 1 0 4807 0 1 9480
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_40
timestamp 1543373569
transform 1 0 4807 0 -1 9480
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_41
timestamp 1543373569
transform 1 0 4807 0 1 8690
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_42
timestamp 1543373569
transform 1 0 4807 0 -1 8690
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_43
timestamp 1543373569
transform 1 0 4807 0 1 7900
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_44
timestamp 1543373569
transform 1 0 4807 0 -1 7900
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_45
timestamp 1543373569
transform 1 0 4807 0 1 7110
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_46
timestamp 1543373569
transform 1 0 4807 0 -1 7110
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_47
timestamp 1543373569
transform 1 0 4807 0 1 6320
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_48
timestamp 1543373569
transform 1 0 4807 0 -1 6320
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_49
timestamp 1543373569
transform 1 0 4807 0 1 5530
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_50
timestamp 1543373569
transform 1 0 4807 0 -1 5530
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_51
timestamp 1543373569
transform 1 0 4807 0 1 4740
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_52
timestamp 1543373569
transform 1 0 4807 0 -1 4740
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_53
timestamp 1543373569
transform 1 0 4807 0 1 3950
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_54
timestamp 1543373569
transform 1 0 4807 0 -1 3950
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_55
timestamp 1543373569
transform 1 0 4807 0 1 3160
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_56
timestamp 1543373569
transform 1 0 4807 0 -1 3160
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_57
timestamp 1543373569
transform 1 0 4807 0 1 2370
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_58
timestamp 1543373569
transform 1 0 4807 0 -1 2370
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_59
timestamp 1543373569
transform 1 0 4807 0 1 1580
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_60
timestamp 1543373569
transform 1 0 4807 0 -1 1580
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_61
timestamp 1543373569
transform 1 0 4807 0 1 790
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_62
timestamp 1543373569
transform 1 0 4807 0 -1 790
box 0 -60 2072 490
use subbyte2_and3_dec  subbyte2_and3_dec_63
timestamp 1543373569
transform 1 0 4807 0 1 0
box 0 -60 2072 490
use subbyte2_hierarchical_predecode2x4  subbyte2_hierarchical_predecode2x4_0
timestamp 1543373569
transform 1 0 527 0 1 4740
box 61 -56 3178 1636
use subbyte2_hierarchical_predecode2x4  subbyte2_hierarchical_predecode2x4_1
timestamp 1543373569
transform 1 0 527 0 1 2370
box 61 -56 3178 1636
use subbyte2_hierarchical_predecode2x4  subbyte2_hierarchical_predecode2x4_2
timestamp 1543373569
transform 1 0 527 0 1 0
box 61 -56 3178 1636
<< labels >>
rlabel metal1 s 19 0 47 6320 4 addr_0
port 3 nsew
rlabel metal1 s 99 0 127 6320 4 addr_1
port 5 nsew
rlabel metal1 s 179 0 207 6320 4 addr_2
port 7 nsew
rlabel metal1 s 259 0 287 6320 4 addr_3
port 9 nsew
rlabel metal1 s 339 0 367 6320 4 addr_4
port 11 nsew
rlabel metal1 s 419 0 447 6320 4 addr_5
port 13 nsew
rlabel locali s 6572 120 6572 120 4 decode_0
port 14 nsew
rlabel locali s 6572 670 6572 670 4 decode_1
port 15 nsew
rlabel locali s 6572 910 6572 910 4 decode_2
port 16 nsew
rlabel locali s 6572 1460 6572 1460 4 decode_3
port 17 nsew
rlabel locali s 6572 1700 6572 1700 4 decode_4
port 18 nsew
rlabel locali s 6572 2250 6572 2250 4 decode_5
port 19 nsew
rlabel locali s 6572 2490 6572 2490 4 decode_6
port 20 nsew
rlabel locali s 6572 3040 6572 3040 4 decode_7
port 21 nsew
rlabel locali s 6572 3280 6572 3280 4 decode_8
port 22 nsew
rlabel locali s 6572 3830 6572 3830 4 decode_9
port 23 nsew
rlabel locali s 6572 4070 6572 4070 4 decode_10
port 24 nsew
rlabel locali s 6572 4620 6572 4620 4 decode_11
port 25 nsew
rlabel locali s 6572 4860 6572 4860 4 decode_12
port 26 nsew
rlabel locali s 6572 5410 6572 5410 4 decode_13
port 27 nsew
rlabel locali s 6572 5650 6572 5650 4 decode_14
port 28 nsew
rlabel locali s 6572 6200 6572 6200 4 decode_15
port 29 nsew
rlabel locali s 6572 6440 6572 6440 4 decode_16
port 30 nsew
rlabel locali s 6572 6990 6572 6990 4 decode_17
port 31 nsew
rlabel locali s 6572 7230 6572 7230 4 decode_18
port 32 nsew
rlabel locali s 6572 7780 6572 7780 4 decode_19
port 33 nsew
rlabel locali s 6572 8020 6572 8020 4 decode_20
port 34 nsew
rlabel locali s 6572 8570 6572 8570 4 decode_21
port 35 nsew
rlabel locali s 6572 8810 6572 8810 4 decode_22
port 36 nsew
rlabel locali s 6572 9360 6572 9360 4 decode_23
port 37 nsew
rlabel locali s 6572 9600 6572 9600 4 decode_24
port 38 nsew
rlabel locali s 6572 10150 6572 10150 4 decode_25
port 39 nsew
rlabel locali s 6572 10390 6572 10390 4 decode_26
port 40 nsew
rlabel locali s 6572 10940 6572 10940 4 decode_27
port 41 nsew
rlabel locali s 6572 11180 6572 11180 4 decode_28
port 42 nsew
rlabel locali s 6572 11730 6572 11730 4 decode_29
port 43 nsew
rlabel locali s 6572 11970 6572 11970 4 decode_30
port 44 nsew
rlabel locali s 6572 12520 6572 12520 4 decode_31
port 45 nsew
rlabel locali s 6572 12760 6572 12760 4 decode_32
port 46 nsew
rlabel locali s 6572 13310 6572 13310 4 decode_33
port 47 nsew
rlabel locali s 6572 13550 6572 13550 4 decode_34
port 48 nsew
rlabel locali s 6572 14100 6572 14100 4 decode_35
port 49 nsew
rlabel locali s 6572 14340 6572 14340 4 decode_36
port 50 nsew
rlabel locali s 6572 14890 6572 14890 4 decode_37
port 51 nsew
rlabel locali s 6572 15130 6572 15130 4 decode_38
port 52 nsew
rlabel locali s 6572 15680 6572 15680 4 decode_39
port 53 nsew
rlabel locali s 6572 15920 6572 15920 4 decode_40
port 54 nsew
rlabel locali s 6572 16470 6572 16470 4 decode_41
port 55 nsew
rlabel locali s 6572 16710 6572 16710 4 decode_42
port 56 nsew
rlabel locali s 6572 17260 6572 17260 4 decode_43
port 57 nsew
rlabel locali s 6572 17500 6572 17500 4 decode_44
port 58 nsew
rlabel locali s 6572 18050 6572 18050 4 decode_45
port 59 nsew
rlabel locali s 6572 18290 6572 18290 4 decode_46
port 60 nsew
rlabel locali s 6572 18840 6572 18840 4 decode_47
port 61 nsew
rlabel locali s 6572 19080 6572 19080 4 decode_48
port 62 nsew
rlabel locali s 6572 19630 6572 19630 4 decode_49
port 63 nsew
rlabel locali s 6572 19870 6572 19870 4 decode_50
port 64 nsew
rlabel locali s 6572 20420 6572 20420 4 decode_51
port 65 nsew
rlabel locali s 6572 20660 6572 20660 4 decode_52
port 66 nsew
rlabel locali s 6572 21210 6572 21210 4 decode_53
port 67 nsew
rlabel locali s 6572 21450 6572 21450 4 decode_54
port 68 nsew
rlabel locali s 6572 22000 6572 22000 4 decode_55
port 69 nsew
rlabel locali s 6572 22240 6572 22240 4 decode_56
port 70 nsew
rlabel locali s 6572 22790 6572 22790 4 decode_57
port 71 nsew
rlabel locali s 6572 23030 6572 23030 4 decode_58
port 72 nsew
rlabel locali s 6572 23580 6572 23580 4 decode_59
port 73 nsew
rlabel locali s 6572 23820 6572 23820 4 decode_60
port 74 nsew
rlabel locali s 6572 24370 6572 24370 4 decode_61
port 75 nsew
rlabel locali s 6572 24610 6572 24610 4 decode_62
port 76 nsew
rlabel locali s 6572 25160 6572 25160 4 decode_63
port 77 nsew
rlabel metal3 s 3490 346 3588 444 4 vdd
port 79 nsew
rlabel metal3 s 3490 1136 3588 1234 4 vdd
port 79 nsew
rlabel metal4 s 6694 -33 6760 25341 4 vdd
port 79 nsew
rlabel metal4 s 5494 -33 5560 25341 4 vdd
port 79 nsew
rlabel metal3 s 2715 353 2813 451 4 vdd
port 79 nsew
rlabel metal3 s 3490 5876 3588 5974 4 vdd
port 79 nsew
rlabel metal3 s 2715 5093 2813 5191 4 vdd
port 79 nsew
rlabel metal3 s 2715 1143 2813 1241 4 vdd
port 79 nsew
rlabel metal3 s 1392 2716 1490 2814 4 vdd
port 79 nsew
rlabel metal3 s 2715 2723 2813 2821 4 vdd
port 79 nsew
rlabel metal3 s 1392 346 1490 444 4 vdd
port 79 nsew
rlabel metal3 s 1392 5086 1490 5184 4 vdd
port 79 nsew
rlabel metal3 s 3490 5086 3588 5184 4 vdd
port 79 nsew
rlabel metal3 s 2715 3513 2813 3611 4 vdd
port 79 nsew
rlabel metal3 s 2715 5883 2813 5981 4 vdd
port 79 nsew
rlabel metal3 s 3490 2716 3588 2814 4 vdd
port 79 nsew
rlabel metal4 s 5926 -33 5992 25341 4 vdd
port 79 nsew
rlabel metal3 s 3490 3506 3588 3604 4 vdd
port 79 nsew
rlabel metal3 s 3094 5876 3192 5974 4 gnd
port 81 nsew
rlabel metal3 s 3094 2716 3192 2814 4 gnd
port 81 nsew
rlabel metal3 s 2290 5883 2388 5981 4 gnd
port 81 nsew
rlabel metal3 s 3094 1136 3192 1234 4 gnd
port 81 nsew
rlabel metal3 s 3094 5086 3192 5184 4 gnd
port 81 nsew
rlabel metal4 s 6270 -33 6336 25341 4 gnd
port 81 nsew
rlabel metal3 s 996 346 1094 444 4 gnd
port 81 nsew
rlabel metal3 s 2290 353 2388 451 4 gnd
port 81 nsew
rlabel metal3 s 3094 346 3192 444 4 gnd
port 81 nsew
rlabel metal3 s 2290 3513 2388 3611 4 gnd
port 81 nsew
rlabel metal3 s 996 5086 1094 5184 4 gnd
port 81 nsew
rlabel metal3 s 996 2716 1094 2814 4 gnd
port 81 nsew
rlabel metal3 s 2290 2723 2388 2821 4 gnd
port 81 nsew
rlabel metal3 s 3094 3506 3192 3604 4 gnd
port 81 nsew
rlabel metal3 s 2290 1143 2388 1241 4 gnd
port 81 nsew
rlabel metal4 s 5022 -33 5088 25341 4 gnd
port 81 nsew
rlabel metal3 s 2290 5093 2388 5191 4 gnd
port 81 nsew
<< properties >>
string FIXED_BBOX 0 0 6861 25308
<< end >>
