magic
tech sky130A
magscale 1 2
timestamp 1543373562
<< checkpaint >>
rect -1260 -1260 47072 43184
<< locali >>
rect 39395 41188 39429 41204
rect 39395 41138 39429 41154
rect 39395 39698 39429 39714
rect 39395 39648 39429 39664
rect 39395 38360 39429 38376
rect 39395 38310 39429 38326
rect 39395 36870 39429 36886
rect 39395 36820 39429 36836
rect 34877 33763 34911 33779
rect 34911 33729 35057 33763
rect 34877 33713 34911 33729
rect 10817 33523 10851 33539
rect 10677 33489 10817 33523
rect 10817 33473 10851 33489
rect 34877 33523 34911 33539
rect 34911 33489 35051 33523
rect 34877 33473 34911 33489
rect 10817 32973 10851 32989
rect 10677 32939 10817 32973
rect 10817 32923 10851 32939
rect 34877 32973 34911 32989
rect 34911 32939 35051 32973
rect 34877 32923 34911 32939
rect 10817 32733 10851 32749
rect 10677 32699 10817 32733
rect 10817 32683 10851 32699
rect 34877 32733 34911 32749
rect 34911 32699 35051 32733
rect 34877 32683 34911 32699
rect 10817 32183 10851 32199
rect 10677 32149 10817 32183
rect 10817 32133 10851 32149
rect 34877 32183 34911 32199
rect 34911 32149 35051 32183
rect 34877 32133 34911 32149
rect 10817 31943 10851 31959
rect 10677 31909 10817 31943
rect 10817 31893 10851 31909
rect 34877 31943 34911 31959
rect 34911 31909 35051 31943
rect 34877 31893 34911 31909
rect 10817 31393 10851 31409
rect 10677 31359 10817 31393
rect 10817 31343 10851 31359
rect 34877 31393 34911 31409
rect 34911 31359 35051 31393
rect 34877 31343 34911 31359
rect 10817 31153 10851 31169
rect 10677 31119 10817 31153
rect 10817 31103 10851 31119
rect 34877 31153 34911 31169
rect 34911 31119 35051 31153
rect 34877 31103 34911 31119
rect 10817 30603 10851 30619
rect 10677 30569 10817 30603
rect 10817 30553 10851 30569
rect 34877 30603 34911 30619
rect 34911 30569 35051 30603
rect 34877 30553 34911 30569
rect 10817 30363 10851 30379
rect 10677 30329 10817 30363
rect 10817 30313 10851 30329
rect 34877 30363 34911 30379
rect 34911 30329 35051 30363
rect 34877 30313 34911 30329
rect 10817 29813 10851 29829
rect 10677 29779 10817 29813
rect 10817 29763 10851 29779
rect 34877 29813 34911 29829
rect 34911 29779 35051 29813
rect 34877 29763 34911 29779
rect 10817 29573 10851 29589
rect 10677 29539 10817 29573
rect 10817 29523 10851 29539
rect 34877 29573 34911 29589
rect 34911 29539 35051 29573
rect 34877 29523 34911 29539
rect 10817 29023 10851 29039
rect 10677 28989 10817 29023
rect 10817 28973 10851 28989
rect 34877 29023 34911 29039
rect 34911 28989 35051 29023
rect 34877 28973 34911 28989
rect 10817 28783 10851 28799
rect 10677 28749 10817 28783
rect 10817 28733 10851 28749
rect 34877 28783 34911 28799
rect 34911 28749 35051 28783
rect 34877 28733 34911 28749
rect 10817 28233 10851 28249
rect 10677 28199 10817 28233
rect 10817 28183 10851 28199
rect 34877 28233 34911 28249
rect 34911 28199 35051 28233
rect 34877 28183 34911 28199
rect 10817 27993 10851 28009
rect 10677 27959 10817 27993
rect 10817 27943 10851 27959
rect 34877 27993 34911 28009
rect 34911 27959 35051 27993
rect 34877 27943 34911 27959
rect 10817 27443 10851 27459
rect 10677 27409 10817 27443
rect 10817 27393 10851 27409
rect 34877 27443 34911 27459
rect 34911 27409 35051 27443
rect 34877 27393 34911 27409
rect 10817 27203 10851 27219
rect 10677 27169 10817 27203
rect 10817 27153 10851 27169
rect 34877 27203 34911 27219
rect 34911 27169 35051 27203
rect 34877 27153 34911 27169
rect 10817 26653 10851 26669
rect 10677 26619 10817 26653
rect 10817 26603 10851 26619
rect 34877 26653 34911 26669
rect 34911 26619 35051 26653
rect 34877 26603 34911 26619
rect 10817 26413 10851 26429
rect 10677 26379 10817 26413
rect 10817 26363 10851 26379
rect 34877 26413 34911 26429
rect 34911 26379 35051 26413
rect 34877 26363 34911 26379
rect 10817 25863 10851 25879
rect 10677 25829 10817 25863
rect 10817 25813 10851 25829
rect 34877 25863 34911 25879
rect 34911 25829 35051 25863
rect 34877 25813 34911 25829
rect 10817 25623 10851 25639
rect 10677 25589 10817 25623
rect 10817 25573 10851 25589
rect 34877 25623 34911 25639
rect 34911 25589 35051 25623
rect 34877 25573 34911 25589
rect 10817 25073 10851 25089
rect 10677 25039 10817 25073
rect 10817 25023 10851 25039
rect 34877 25073 34911 25089
rect 34911 25039 35051 25073
rect 34877 25023 34911 25039
rect 10817 24833 10851 24849
rect 10677 24799 10817 24833
rect 10817 24783 10851 24799
rect 34877 24833 34911 24849
rect 34911 24799 35051 24833
rect 34877 24783 34911 24799
rect 10817 24283 10851 24299
rect 10677 24249 10817 24283
rect 10817 24233 10851 24249
rect 34877 24283 34911 24299
rect 34911 24249 35051 24283
rect 34877 24233 34911 24249
rect 10817 24043 10851 24059
rect 10677 24009 10817 24043
rect 10817 23993 10851 24009
rect 34877 24043 34911 24059
rect 34911 24009 35051 24043
rect 34877 23993 34911 24009
rect 10817 23493 10851 23509
rect 10677 23459 10817 23493
rect 10817 23443 10851 23459
rect 34877 23493 34911 23509
rect 34911 23459 35051 23493
rect 34877 23443 34911 23459
rect 10817 23253 10851 23269
rect 10677 23219 10817 23253
rect 10817 23203 10851 23219
rect 34877 23253 34911 23269
rect 34911 23219 35051 23253
rect 34877 23203 34911 23219
rect 10817 22703 10851 22719
rect 10677 22669 10817 22703
rect 10817 22653 10851 22669
rect 34877 22703 34911 22719
rect 34911 22669 35051 22703
rect 34877 22653 34911 22669
rect 10817 22463 10851 22479
rect 10677 22429 10817 22463
rect 10817 22413 10851 22429
rect 34877 22463 34911 22479
rect 34911 22429 35051 22463
rect 34877 22413 34911 22429
rect 10817 21913 10851 21929
rect 10677 21879 10817 21913
rect 10817 21863 10851 21879
rect 34877 21913 34911 21929
rect 34911 21879 35051 21913
rect 34877 21863 34911 21879
rect 10817 21673 10851 21689
rect 10677 21639 10817 21673
rect 10817 21623 10851 21639
rect 34877 21673 34911 21689
rect 34911 21639 35051 21673
rect 34877 21623 34911 21639
rect 10817 21123 10851 21139
rect 10677 21089 10817 21123
rect 10817 21073 10851 21089
rect 34877 21123 34911 21139
rect 34911 21089 35051 21123
rect 34877 21073 34911 21089
rect 10817 20883 10851 20899
rect 10677 20849 10817 20883
rect 10817 20833 10851 20849
rect 34877 20883 34911 20899
rect 34911 20849 35051 20883
rect 34877 20833 34911 20849
rect 10817 20333 10851 20349
rect 10677 20299 10817 20333
rect 10817 20283 10851 20299
rect 34877 20333 34911 20349
rect 34911 20299 35051 20333
rect 34877 20283 34911 20299
rect 10817 20093 10851 20109
rect 10677 20059 10817 20093
rect 10817 20043 10851 20059
rect 34877 20093 34911 20109
rect 34911 20059 35051 20093
rect 34877 20043 34911 20059
rect 10817 19543 10851 19559
rect 10677 19509 10817 19543
rect 10817 19493 10851 19509
rect 34877 19543 34911 19559
rect 34911 19509 35051 19543
rect 34877 19493 34911 19509
rect 10817 19303 10851 19319
rect 10677 19269 10817 19303
rect 10817 19253 10851 19269
rect 34877 19303 34911 19319
rect 34911 19269 35051 19303
rect 34877 19253 34911 19269
rect 10817 18753 10851 18769
rect 10677 18719 10817 18753
rect 10817 18703 10851 18719
rect 34877 18753 34911 18769
rect 34911 18719 35051 18753
rect 34877 18703 34911 18719
rect 10817 18513 10851 18529
rect 10677 18479 10817 18513
rect 10817 18463 10851 18479
rect 34877 18513 34911 18529
rect 34911 18479 35051 18513
rect 34877 18463 34911 18479
rect 10817 17963 10851 17979
rect 10677 17929 10817 17963
rect 10817 17913 10851 17929
rect 34877 17963 34911 17979
rect 34911 17929 35051 17963
rect 34877 17913 34911 17929
rect 10817 17723 10851 17739
rect 10677 17689 10817 17723
rect 10817 17673 10851 17689
rect 34877 17723 34911 17739
rect 34911 17689 35051 17723
rect 34877 17673 34911 17689
rect 10817 17173 10851 17189
rect 10677 17139 10817 17173
rect 10817 17123 10851 17139
rect 34877 17173 34911 17189
rect 34911 17139 35051 17173
rect 34877 17123 34911 17139
rect 10817 16933 10851 16949
rect 10677 16899 10817 16933
rect 10817 16883 10851 16899
rect 34877 16933 34911 16949
rect 34911 16899 35051 16933
rect 34877 16883 34911 16899
rect 10817 16383 10851 16399
rect 10677 16349 10817 16383
rect 10817 16333 10851 16349
rect 34877 16383 34911 16399
rect 34911 16349 35051 16383
rect 34877 16333 34911 16349
rect 10817 16143 10851 16159
rect 10677 16109 10817 16143
rect 10817 16093 10851 16109
rect 34877 16143 34911 16159
rect 34911 16109 35051 16143
rect 34877 16093 34911 16109
rect 10817 15593 10851 15609
rect 10677 15559 10817 15593
rect 10817 15543 10851 15559
rect 34877 15593 34911 15609
rect 34911 15559 35051 15593
rect 34877 15543 34911 15559
rect 10817 15353 10851 15369
rect 10677 15319 10817 15353
rect 10817 15303 10851 15319
rect 34877 15353 34911 15369
rect 34911 15319 35051 15353
rect 34877 15303 34911 15319
rect 10817 14803 10851 14819
rect 10677 14769 10817 14803
rect 10817 14753 10851 14769
rect 34877 14803 34911 14819
rect 34911 14769 35051 14803
rect 34877 14753 34911 14769
rect 10817 14563 10851 14579
rect 10677 14529 10817 14563
rect 10817 14513 10851 14529
rect 34877 14563 34911 14579
rect 34911 14529 35051 14563
rect 34877 14513 34911 14529
rect 10817 14013 10851 14029
rect 10677 13979 10817 14013
rect 10817 13963 10851 13979
rect 34877 14013 34911 14029
rect 34911 13979 35051 14013
rect 34877 13963 34911 13979
rect 10817 13773 10851 13789
rect 10677 13739 10817 13773
rect 10817 13723 10851 13739
rect 34877 13773 34911 13789
rect 34911 13739 35051 13773
rect 34877 13723 34911 13739
rect 10817 13223 10851 13239
rect 10677 13189 10817 13223
rect 10817 13173 10851 13189
rect 34877 13223 34911 13239
rect 34911 13189 35051 13223
rect 34877 13173 34911 13189
rect 10817 12983 10851 12999
rect 10677 12949 10817 12983
rect 10817 12933 10851 12949
rect 34877 12983 34911 12999
rect 34911 12949 35051 12983
rect 34877 12933 34911 12949
rect 10817 12433 10851 12449
rect 10677 12399 10817 12433
rect 10817 12383 10851 12399
rect 34877 12433 34911 12449
rect 34911 12399 35051 12433
rect 34877 12383 34911 12399
rect 10817 12193 10851 12209
rect 10677 12159 10817 12193
rect 10817 12143 10851 12159
rect 34877 12193 34911 12209
rect 34911 12159 35051 12193
rect 34877 12143 34911 12159
rect 10817 11643 10851 11659
rect 10677 11609 10817 11643
rect 10817 11593 10851 11609
rect 34877 11643 34911 11659
rect 34911 11609 35051 11643
rect 34877 11593 34911 11609
rect 10817 11403 10851 11419
rect 10677 11369 10817 11403
rect 10817 11353 10851 11369
rect 34877 11403 34911 11419
rect 34911 11369 35051 11403
rect 34877 11353 34911 11369
rect 10817 10853 10851 10869
rect 10677 10819 10817 10853
rect 10817 10803 10851 10819
rect 34877 10853 34911 10869
rect 34911 10819 35051 10853
rect 34877 10803 34911 10819
rect 10817 10613 10851 10629
rect 10677 10579 10817 10613
rect 10817 10563 10851 10579
rect 34877 10613 34911 10629
rect 34911 10579 35051 10613
rect 34877 10563 34911 10579
rect 10817 10063 10851 10079
rect 10677 10029 10817 10063
rect 10817 10013 10851 10029
rect 34877 10063 34911 10079
rect 34911 10029 35051 10063
rect 34877 10013 34911 10029
rect 10817 9823 10851 9839
rect 10677 9789 10817 9823
rect 10817 9773 10851 9789
rect 34877 9823 34911 9839
rect 34911 9789 35051 9823
rect 34877 9773 34911 9789
rect 10817 9273 10851 9289
rect 10677 9239 10817 9273
rect 10817 9223 10851 9239
rect 34877 9273 34911 9289
rect 34911 9239 35051 9273
rect 34877 9223 34911 9239
rect 10817 9033 10851 9049
rect 10677 8999 10817 9033
rect 10817 8983 10851 8999
rect 34877 9033 34911 9049
rect 34911 8999 35051 9033
rect 34877 8983 34911 8999
rect 10817 8483 10851 8499
rect 10677 8449 10817 8483
rect 10817 8433 10851 8449
rect 34877 8483 34911 8499
rect 34911 8449 35051 8483
rect 34877 8433 34911 8449
rect 10817 8243 10851 8259
rect 10671 8209 10817 8243
rect 10817 8193 10851 8209
rect 6299 5086 6333 5102
rect 6299 5036 6333 5052
rect 6299 3596 6333 3612
rect 6299 3546 6333 3562
rect 6299 2258 6333 2274
rect 6299 2208 6333 2224
rect 6299 768 6333 784
rect 6299 718 6333 734
<< viali >>
rect 39395 41154 39429 41188
rect 39395 39664 39429 39698
rect 39395 38326 39429 38360
rect 39395 36836 39429 36870
rect 34877 33729 34911 33763
rect 10817 33489 10851 33523
rect 34877 33489 34911 33523
rect 10817 32939 10851 32973
rect 34877 32939 34911 32973
rect 10817 32699 10851 32733
rect 34877 32699 34911 32733
rect 10817 32149 10851 32183
rect 34877 32149 34911 32183
rect 10817 31909 10851 31943
rect 34877 31909 34911 31943
rect 10817 31359 10851 31393
rect 34877 31359 34911 31393
rect 10817 31119 10851 31153
rect 34877 31119 34911 31153
rect 10817 30569 10851 30603
rect 34877 30569 34911 30603
rect 10817 30329 10851 30363
rect 34877 30329 34911 30363
rect 10817 29779 10851 29813
rect 34877 29779 34911 29813
rect 10817 29539 10851 29573
rect 34877 29539 34911 29573
rect 10817 28989 10851 29023
rect 34877 28989 34911 29023
rect 10817 28749 10851 28783
rect 34877 28749 34911 28783
rect 10817 28199 10851 28233
rect 34877 28199 34911 28233
rect 10817 27959 10851 27993
rect 34877 27959 34911 27993
rect 10817 27409 10851 27443
rect 34877 27409 34911 27443
rect 10817 27169 10851 27203
rect 34877 27169 34911 27203
rect 10817 26619 10851 26653
rect 34877 26619 34911 26653
rect 10817 26379 10851 26413
rect 34877 26379 34911 26413
rect 10817 25829 10851 25863
rect 34877 25829 34911 25863
rect 10817 25589 10851 25623
rect 34877 25589 34911 25623
rect 10817 25039 10851 25073
rect 34877 25039 34911 25073
rect 10817 24799 10851 24833
rect 34877 24799 34911 24833
rect 10817 24249 10851 24283
rect 34877 24249 34911 24283
rect 10817 24009 10851 24043
rect 34877 24009 34911 24043
rect 10817 23459 10851 23493
rect 34877 23459 34911 23493
rect 10817 23219 10851 23253
rect 34877 23219 34911 23253
rect 10817 22669 10851 22703
rect 34877 22669 34911 22703
rect 10817 22429 10851 22463
rect 34877 22429 34911 22463
rect 10817 21879 10851 21913
rect 34877 21879 34911 21913
rect 10817 21639 10851 21673
rect 34877 21639 34911 21673
rect 10817 21089 10851 21123
rect 34877 21089 34911 21123
rect 10817 20849 10851 20883
rect 34877 20849 34911 20883
rect 10817 20299 10851 20333
rect 34877 20299 34911 20333
rect 10817 20059 10851 20093
rect 34877 20059 34911 20093
rect 10817 19509 10851 19543
rect 34877 19509 34911 19543
rect 10817 19269 10851 19303
rect 34877 19269 34911 19303
rect 10817 18719 10851 18753
rect 34877 18719 34911 18753
rect 10817 18479 10851 18513
rect 34877 18479 34911 18513
rect 10817 17929 10851 17963
rect 34877 17929 34911 17963
rect 10817 17689 10851 17723
rect 34877 17689 34911 17723
rect 10817 17139 10851 17173
rect 34877 17139 34911 17173
rect 10817 16899 10851 16933
rect 34877 16899 34911 16933
rect 10817 16349 10851 16383
rect 34877 16349 34911 16383
rect 10817 16109 10851 16143
rect 34877 16109 34911 16143
rect 10817 15559 10851 15593
rect 34877 15559 34911 15593
rect 10817 15319 10851 15353
rect 34877 15319 34911 15353
rect 10817 14769 10851 14803
rect 34877 14769 34911 14803
rect 10817 14529 10851 14563
rect 34877 14529 34911 14563
rect 10817 13979 10851 14013
rect 34877 13979 34911 14013
rect 10817 13739 10851 13773
rect 34877 13739 34911 13773
rect 10817 13189 10851 13223
rect 34877 13189 34911 13223
rect 10817 12949 10851 12983
rect 34877 12949 34911 12983
rect 10817 12399 10851 12433
rect 34877 12399 34911 12433
rect 10817 12159 10851 12193
rect 34877 12159 34911 12193
rect 10817 11609 10851 11643
rect 34877 11609 34911 11643
rect 10817 11369 10851 11403
rect 34877 11369 34911 11403
rect 10817 10819 10851 10853
rect 34877 10819 34911 10853
rect 10817 10579 10851 10613
rect 34877 10579 34911 10613
rect 10817 10029 10851 10063
rect 34877 10029 34911 10063
rect 10817 9789 10851 9823
rect 34877 9789 34911 9823
rect 10817 9239 10851 9273
rect 34877 9239 34911 9273
rect 10817 8999 10851 9033
rect 34877 8999 34911 9033
rect 10817 8449 10851 8483
rect 34877 8449 34911 8483
rect 10817 8209 10851 8243
rect 6299 5052 6333 5086
rect 6299 3562 6333 3596
rect 6299 2224 6333 2258
rect 6299 734 6333 768
<< metal1 >>
rect 39380 41145 39386 41197
rect 39438 41145 39444 41197
rect 41450 41142 41496 41200
rect 12984 40484 13030 40634
rect 15480 40484 15526 40634
rect 17976 40484 18022 40634
rect 20472 40484 20518 40634
rect 22968 40484 23014 40634
rect 25464 40484 25510 40634
rect 27960 40484 28006 40634
rect 30456 40484 30502 40634
rect 39380 39655 39386 39707
rect 39438 39655 39444 39707
rect 41326 39652 41372 39710
rect 39380 38317 39386 38369
rect 39438 38317 39444 38369
rect 39380 36827 39386 36879
rect 39438 36827 39444 36879
rect 32896 35488 32902 35540
rect 32954 35488 32960 35540
rect 32914 35390 32942 35488
rect 12946 34556 12974 34668
rect 13410 34556 13438 34668
rect 12946 34528 13206 34556
rect 13178 34416 13206 34528
rect 13250 34528 13438 34556
rect 13570 34556 13598 34668
rect 14034 34556 14062 34668
rect 13570 34528 13758 34556
rect 13250 34416 13278 34528
rect 13730 34416 13758 34528
rect 13802 34528 14062 34556
rect 14194 34556 14222 34668
rect 14658 34556 14686 34668
rect 14194 34528 14454 34556
rect 13802 34416 13830 34528
rect 14426 34416 14454 34528
rect 14498 34528 14686 34556
rect 14818 34556 14846 34668
rect 15282 34556 15310 34668
rect 14818 34528 15006 34556
rect 14498 34416 14526 34528
rect 14978 34416 15006 34528
rect 15050 34528 15310 34556
rect 15442 34556 15470 34668
rect 15906 34556 15934 34668
rect 15442 34528 15702 34556
rect 15050 34416 15078 34528
rect 15674 34416 15702 34528
rect 15746 34528 15934 34556
rect 16066 34556 16094 34668
rect 16530 34556 16558 34668
rect 16066 34528 16254 34556
rect 15746 34416 15774 34528
rect 16226 34416 16254 34528
rect 16298 34528 16558 34556
rect 16690 34556 16718 34668
rect 17154 34556 17182 34668
rect 16690 34528 16950 34556
rect 16298 34416 16326 34528
rect 16922 34416 16950 34528
rect 16994 34528 17182 34556
rect 17314 34556 17342 34668
rect 17778 34556 17806 34668
rect 17314 34528 17502 34556
rect 16994 34416 17022 34528
rect 17474 34416 17502 34528
rect 17546 34528 17806 34556
rect 17938 34556 17966 34668
rect 18402 34556 18430 34668
rect 17938 34528 18198 34556
rect 17546 34416 17574 34528
rect 18170 34416 18198 34528
rect 18242 34528 18430 34556
rect 18562 34556 18590 34668
rect 19026 34556 19054 34668
rect 18562 34528 18750 34556
rect 18242 34416 18270 34528
rect 18722 34416 18750 34528
rect 18794 34528 19054 34556
rect 19186 34556 19214 34668
rect 19650 34556 19678 34668
rect 19186 34528 19446 34556
rect 18794 34416 18822 34528
rect 19418 34416 19446 34528
rect 19490 34528 19678 34556
rect 19810 34556 19838 34668
rect 20274 34556 20302 34668
rect 19810 34528 19998 34556
rect 19490 34416 19518 34528
rect 19970 34416 19998 34528
rect 20042 34528 20302 34556
rect 20434 34556 20462 34668
rect 20898 34556 20926 34668
rect 20434 34528 20694 34556
rect 20042 34416 20070 34528
rect 20666 34416 20694 34528
rect 20738 34528 20926 34556
rect 21058 34556 21086 34668
rect 21522 34556 21550 34668
rect 21058 34528 21246 34556
rect 20738 34416 20766 34528
rect 21218 34416 21246 34528
rect 21290 34528 21550 34556
rect 21682 34556 21710 34668
rect 22146 34556 22174 34668
rect 21682 34528 21942 34556
rect 21290 34416 21318 34528
rect 21914 34416 21942 34528
rect 21986 34528 22174 34556
rect 22306 34556 22334 34668
rect 22770 34556 22798 34668
rect 22306 34528 22494 34556
rect 21986 34416 22014 34528
rect 22466 34416 22494 34528
rect 22538 34528 22798 34556
rect 22930 34556 22958 34668
rect 23394 34556 23422 34668
rect 22930 34528 23190 34556
rect 22538 34416 22566 34528
rect 23162 34416 23190 34528
rect 23234 34528 23422 34556
rect 23554 34556 23582 34668
rect 24018 34556 24046 34668
rect 23554 34528 23742 34556
rect 23234 34416 23262 34528
rect 23714 34416 23742 34528
rect 23786 34528 24046 34556
rect 24178 34556 24206 34668
rect 24642 34556 24670 34668
rect 24178 34528 24438 34556
rect 23786 34416 23814 34528
rect 24410 34416 24438 34528
rect 24482 34528 24670 34556
rect 24802 34556 24830 34668
rect 25266 34556 25294 34668
rect 24802 34528 24990 34556
rect 24482 34416 24510 34528
rect 24962 34416 24990 34528
rect 25034 34528 25294 34556
rect 25426 34556 25454 34668
rect 25890 34556 25918 34668
rect 25426 34528 25686 34556
rect 25034 34416 25062 34528
rect 25658 34416 25686 34528
rect 25730 34528 25918 34556
rect 26050 34556 26078 34668
rect 26514 34556 26542 34668
rect 26050 34528 26238 34556
rect 25730 34416 25758 34528
rect 26210 34416 26238 34528
rect 26282 34528 26542 34556
rect 26674 34556 26702 34668
rect 27138 34556 27166 34668
rect 26674 34528 26934 34556
rect 26282 34416 26310 34528
rect 26906 34416 26934 34528
rect 26978 34528 27166 34556
rect 27298 34556 27326 34668
rect 27762 34556 27790 34668
rect 27298 34528 27486 34556
rect 26978 34416 27006 34528
rect 27458 34416 27486 34528
rect 27530 34528 27790 34556
rect 27922 34556 27950 34668
rect 28386 34556 28414 34668
rect 27922 34528 28182 34556
rect 27530 34416 27558 34528
rect 28154 34416 28182 34528
rect 28226 34528 28414 34556
rect 28546 34556 28574 34668
rect 29010 34556 29038 34668
rect 28546 34528 28734 34556
rect 28226 34416 28254 34528
rect 28706 34416 28734 34528
rect 28778 34528 29038 34556
rect 29170 34556 29198 34668
rect 29634 34556 29662 34668
rect 29170 34528 29430 34556
rect 28778 34416 28806 34528
rect 29402 34416 29430 34528
rect 29474 34528 29662 34556
rect 29794 34556 29822 34668
rect 30258 34556 30286 34668
rect 29794 34528 29982 34556
rect 29474 34416 29502 34528
rect 29954 34416 29982 34528
rect 30026 34528 30286 34556
rect 30418 34556 30446 34668
rect 30882 34556 30910 34668
rect 30418 34528 30678 34556
rect 30026 34416 30054 34528
rect 30650 34416 30678 34528
rect 30722 34528 30910 34556
rect 31042 34556 31070 34668
rect 31506 34556 31534 34668
rect 31042 34528 31230 34556
rect 30722 34416 30750 34528
rect 31202 34416 31230 34528
rect 31274 34528 31534 34556
rect 31666 34556 31694 34668
rect 32130 34556 32158 34668
rect 31666 34528 31926 34556
rect 31274 34416 31302 34528
rect 31898 34416 31926 34528
rect 31970 34528 32158 34556
rect 32290 34556 32318 34668
rect 32754 34556 32782 34668
rect 32290 34528 32478 34556
rect 31970 34416 31998 34528
rect 32450 34416 32478 34528
rect 32522 34528 32782 34556
rect 32914 34556 32942 34668
rect 33378 34556 33406 34668
rect 32914 34528 33174 34556
rect 32522 34416 32550 34528
rect 33146 34416 33174 34528
rect 33218 34528 33406 34556
rect 33218 34416 33246 34528
rect 34862 33720 34868 33772
rect 34920 33720 34926 33772
rect 35779 33626 35807 34021
rect 37659 33594 37709 34028
rect 10802 33480 10808 33532
rect 10860 33480 10866 33532
rect 34862 33480 34868 33532
rect 34920 33480 34926 33532
rect 10802 32930 10808 32982
rect 10860 32930 10866 32982
rect 34862 32930 34868 32982
rect 34920 32930 34926 32982
rect 10802 32690 10808 32742
rect 10860 32690 10866 32742
rect 34862 32690 34868 32742
rect 34920 32690 34926 32742
rect 10802 32140 10808 32192
rect 10860 32140 10866 32192
rect 34862 32140 34868 32192
rect 34920 32140 34926 32192
rect 10802 31900 10808 31952
rect 10860 31900 10866 31952
rect 34862 31900 34868 31952
rect 34920 31900 34926 31952
rect 10802 31350 10808 31402
rect 10860 31350 10866 31402
rect 34862 31350 34868 31402
rect 34920 31350 34926 31402
rect 10802 31110 10808 31162
rect 10860 31110 10866 31162
rect 34862 31110 34868 31162
rect 34920 31110 34926 31162
rect 10802 30560 10808 30612
rect 10860 30560 10866 30612
rect 34862 30560 34868 30612
rect 34920 30560 34926 30612
rect 10802 30320 10808 30372
rect 10860 30320 10866 30372
rect 34862 30320 34868 30372
rect 34920 30320 34926 30372
rect 10802 29770 10808 29822
rect 10860 29770 10866 29822
rect 34862 29770 34868 29822
rect 34920 29770 34926 29822
rect 10802 29530 10808 29582
rect 10860 29530 10866 29582
rect 34862 29530 34868 29582
rect 34920 29530 34926 29582
rect 10802 28980 10808 29032
rect 10860 28980 10866 29032
rect 34862 28980 34868 29032
rect 34920 28980 34926 29032
rect 10802 28740 10808 28792
rect 10860 28740 10866 28792
rect 34862 28740 34868 28792
rect 34920 28740 34926 28792
rect 10802 28190 10808 28242
rect 10860 28190 10866 28242
rect 34862 28190 34868 28242
rect 34920 28190 34926 28242
rect 10802 27950 10808 28002
rect 10860 27950 10866 28002
rect 34862 27950 34868 28002
rect 34920 27950 34926 28002
rect 10802 27400 10808 27452
rect 10860 27400 10866 27452
rect 34862 27400 34868 27452
rect 34920 27400 34926 27452
rect 10802 27160 10808 27212
rect 10860 27160 10866 27212
rect 34862 27160 34868 27212
rect 34920 27160 34926 27212
rect 10802 26610 10808 26662
rect 10860 26610 10866 26662
rect 34862 26610 34868 26662
rect 34920 26610 34926 26662
rect 10802 26370 10808 26422
rect 10860 26370 10866 26422
rect 34862 26370 34868 26422
rect 34920 26370 34926 26422
rect 10802 25820 10808 25872
rect 10860 25820 10866 25872
rect 34862 25820 34868 25872
rect 34920 25820 34926 25872
rect 10802 25580 10808 25632
rect 10860 25580 10866 25632
rect 34862 25580 34868 25632
rect 34920 25580 34926 25632
rect 10802 25030 10808 25082
rect 10860 25030 10866 25082
rect 34862 25030 34868 25082
rect 34920 25030 34926 25082
rect 10802 24790 10808 24842
rect 10860 24790 10866 24842
rect 34862 24790 34868 24842
rect 34920 24790 34926 24842
rect 10802 24240 10808 24292
rect 10860 24240 10866 24292
rect 34862 24240 34868 24292
rect 34920 24240 34926 24292
rect 10802 24000 10808 24052
rect 10860 24000 10866 24052
rect 34862 24000 34868 24052
rect 34920 24000 34926 24052
rect 10802 23450 10808 23502
rect 10860 23450 10866 23502
rect 34862 23450 34868 23502
rect 34920 23450 34926 23502
rect 10802 23210 10808 23262
rect 10860 23210 10866 23262
rect 34862 23210 34868 23262
rect 34920 23210 34926 23262
rect 10802 22660 10808 22712
rect 10860 22660 10866 22712
rect 34862 22660 34868 22712
rect 34920 22660 34926 22712
rect 10802 22420 10808 22472
rect 10860 22420 10866 22472
rect 34862 22420 34868 22472
rect 34920 22420 34926 22472
rect 10802 21870 10808 21922
rect 10860 21870 10866 21922
rect 34862 21870 34868 21922
rect 34920 21870 34926 21922
rect 10802 21630 10808 21682
rect 10860 21630 10866 21682
rect 34862 21630 34868 21682
rect 34920 21630 34926 21682
rect 10802 21080 10808 21132
rect 10860 21080 10866 21132
rect 34862 21080 34868 21132
rect 34920 21080 34926 21132
rect 10802 20840 10808 20892
rect 10860 20840 10866 20892
rect 34862 20840 34868 20892
rect 34920 20840 34926 20892
rect 10802 20290 10808 20342
rect 10860 20290 10866 20342
rect 34862 20290 34868 20342
rect 34920 20290 34926 20342
rect 10802 20050 10808 20102
rect 10860 20050 10866 20102
rect 34862 20050 34868 20102
rect 34920 20050 34926 20102
rect 10802 19500 10808 19552
rect 10860 19500 10866 19552
rect 34862 19500 34868 19552
rect 34920 19500 34926 19552
rect 10802 19260 10808 19312
rect 10860 19260 10866 19312
rect 34862 19260 34868 19312
rect 34920 19260 34926 19312
rect 10802 18710 10808 18762
rect 10860 18710 10866 18762
rect 34862 18710 34868 18762
rect 34920 18710 34926 18762
rect 10802 18470 10808 18522
rect 10860 18470 10866 18522
rect 34862 18470 34868 18522
rect 34920 18470 34926 18522
rect 10802 17920 10808 17972
rect 10860 17920 10866 17972
rect 34862 17920 34868 17972
rect 34920 17920 34926 17972
rect 10802 17680 10808 17732
rect 10860 17680 10866 17732
rect 34862 17680 34868 17732
rect 34920 17680 34926 17732
rect 10802 17130 10808 17182
rect 10860 17130 10866 17182
rect 34862 17130 34868 17182
rect 34920 17130 34926 17182
rect 10802 16890 10808 16942
rect 10860 16890 10866 16942
rect 34862 16890 34868 16942
rect 34920 16890 34926 16942
rect 10802 16340 10808 16392
rect 10860 16340 10866 16392
rect 34862 16340 34868 16392
rect 34920 16340 34926 16392
rect 10802 16100 10808 16152
rect 10860 16100 10866 16152
rect 34862 16100 34868 16152
rect 34920 16100 34926 16152
rect 10802 15550 10808 15602
rect 10860 15550 10866 15602
rect 34862 15550 34868 15602
rect 34920 15550 34926 15602
rect 10802 15310 10808 15362
rect 10860 15310 10866 15362
rect 34862 15310 34868 15362
rect 34920 15310 34926 15362
rect 10802 14760 10808 14812
rect 10860 14760 10866 14812
rect 34862 14760 34868 14812
rect 34920 14760 34926 14812
rect 19 8346 47 14666
rect 99 8346 127 14666
rect 179 8346 207 14666
rect 259 8346 287 14666
rect 339 8346 367 14666
rect 419 8346 447 14666
rect 10802 14520 10808 14572
rect 10860 14520 10866 14572
rect 34862 14520 34868 14572
rect 34920 14520 34926 14572
rect 10802 13970 10808 14022
rect 10860 13970 10866 14022
rect 34862 13970 34868 14022
rect 34920 13970 34926 14022
rect 10802 13730 10808 13782
rect 10860 13730 10866 13782
rect 34862 13730 34868 13782
rect 34920 13730 34926 13782
rect 10802 13180 10808 13232
rect 10860 13180 10866 13232
rect 34862 13180 34868 13232
rect 34920 13180 34926 13232
rect 10802 12940 10808 12992
rect 10860 12940 10866 12992
rect 34862 12940 34868 12992
rect 34920 12940 34926 12992
rect 10802 12390 10808 12442
rect 10860 12390 10866 12442
rect 34862 12390 34868 12442
rect 34920 12390 34926 12442
rect 10802 12150 10808 12202
rect 10860 12150 10866 12202
rect 34862 12150 34868 12202
rect 34920 12150 34926 12202
rect 10802 11600 10808 11652
rect 10860 11600 10866 11652
rect 34862 11600 34868 11652
rect 34920 11600 34926 11652
rect 10802 11360 10808 11412
rect 10860 11360 10866 11412
rect 34862 11360 34868 11412
rect 34920 11360 34926 11412
rect 10802 10810 10808 10862
rect 10860 10810 10866 10862
rect 34862 10810 34868 10862
rect 34920 10810 34926 10862
rect 10802 10570 10808 10622
rect 10860 10570 10866 10622
rect 34862 10570 34868 10622
rect 34920 10570 34926 10622
rect 10802 10020 10808 10072
rect 10860 10020 10866 10072
rect 34862 10020 34868 10072
rect 34920 10020 34926 10072
rect 10802 9780 10808 9832
rect 10860 9780 10866 9832
rect 34862 9780 34868 9832
rect 34920 9780 34926 9832
rect 10802 9230 10808 9282
rect 10860 9230 10866 9282
rect 34862 9230 34868 9282
rect 34920 9230 34926 9282
rect 10802 8990 10808 9042
rect 10860 8990 10866 9042
rect 34862 8990 34868 9042
rect 34920 8990 34926 9042
rect 10802 8440 10808 8492
rect 10860 8440 10866 8492
rect 34862 8440 34868 8492
rect 34920 8440 34926 8492
rect 8019 7944 8069 8378
rect 45281 8346 45309 14666
rect 45361 8346 45389 14666
rect 45441 8346 45469 14666
rect 45521 8346 45549 14666
rect 45601 8346 45629 14666
rect 45681 8346 45709 14666
rect 9921 7951 9949 8346
rect 10802 8200 10808 8252
rect 10860 8200 10866 8252
rect 12698 7394 12726 7506
rect 12322 7366 12726 7394
rect 12770 7394 12798 7506
rect 12962 7394 12990 7506
rect 12770 7366 12814 7394
rect 12322 7254 12350 7366
rect 12786 7254 12814 7366
rect 12946 7366 12990 7394
rect 13034 7394 13062 7506
rect 13946 7394 13974 7506
rect 13034 7366 13438 7394
rect 12946 7254 12974 7366
rect 13410 7254 13438 7366
rect 13570 7366 13974 7394
rect 14018 7394 14046 7506
rect 14210 7394 14238 7506
rect 14018 7366 14062 7394
rect 13570 7254 13598 7366
rect 14034 7254 14062 7366
rect 14194 7366 14238 7394
rect 14282 7394 14310 7506
rect 15194 7394 15222 7506
rect 14282 7366 14686 7394
rect 14194 7254 14222 7366
rect 14658 7254 14686 7366
rect 14818 7366 15222 7394
rect 15266 7394 15294 7506
rect 15458 7394 15486 7506
rect 15266 7366 15310 7394
rect 14818 7254 14846 7366
rect 15282 7254 15310 7366
rect 15442 7366 15486 7394
rect 15530 7394 15558 7506
rect 16442 7394 16470 7506
rect 15530 7366 15934 7394
rect 15442 7254 15470 7366
rect 15906 7254 15934 7366
rect 16066 7366 16470 7394
rect 16514 7394 16542 7506
rect 16706 7394 16734 7506
rect 16514 7366 16558 7394
rect 16066 7254 16094 7366
rect 16530 7254 16558 7366
rect 16690 7366 16734 7394
rect 16778 7394 16806 7506
rect 17690 7394 17718 7506
rect 16778 7366 17182 7394
rect 16690 7254 16718 7366
rect 17154 7254 17182 7366
rect 17314 7366 17718 7394
rect 17762 7394 17790 7506
rect 17954 7394 17982 7506
rect 17762 7366 17806 7394
rect 17314 7254 17342 7366
rect 17778 7254 17806 7366
rect 17938 7366 17982 7394
rect 18026 7394 18054 7506
rect 18938 7394 18966 7506
rect 18026 7366 18430 7394
rect 17938 7254 17966 7366
rect 18402 7254 18430 7366
rect 18562 7366 18966 7394
rect 19010 7394 19038 7506
rect 19202 7394 19230 7506
rect 19010 7366 19054 7394
rect 18562 7254 18590 7366
rect 19026 7254 19054 7366
rect 19186 7366 19230 7394
rect 19274 7394 19302 7506
rect 20186 7394 20214 7506
rect 19274 7366 19678 7394
rect 19186 7254 19214 7366
rect 19650 7254 19678 7366
rect 19810 7366 20214 7394
rect 20258 7394 20286 7506
rect 20450 7394 20478 7506
rect 20258 7366 20302 7394
rect 19810 7254 19838 7366
rect 20274 7254 20302 7366
rect 20434 7366 20478 7394
rect 20522 7394 20550 7506
rect 21434 7394 21462 7506
rect 20522 7366 20926 7394
rect 20434 7254 20462 7366
rect 20898 7254 20926 7366
rect 21058 7366 21462 7394
rect 21506 7394 21534 7506
rect 21698 7394 21726 7506
rect 21506 7366 21550 7394
rect 21058 7254 21086 7366
rect 21522 7254 21550 7366
rect 21682 7366 21726 7394
rect 21770 7394 21798 7506
rect 22682 7394 22710 7506
rect 21770 7366 22174 7394
rect 21682 7254 21710 7366
rect 22146 7254 22174 7366
rect 22306 7366 22710 7394
rect 22754 7394 22782 7506
rect 22946 7394 22974 7506
rect 22754 7366 22798 7394
rect 22306 7254 22334 7366
rect 22770 7254 22798 7366
rect 22930 7366 22974 7394
rect 23018 7394 23046 7506
rect 23930 7394 23958 7506
rect 23018 7366 23422 7394
rect 22930 7254 22958 7366
rect 23394 7254 23422 7366
rect 23554 7366 23958 7394
rect 24002 7394 24030 7506
rect 24194 7394 24222 7506
rect 24002 7366 24046 7394
rect 23554 7254 23582 7366
rect 24018 7254 24046 7366
rect 24178 7366 24222 7394
rect 24266 7394 24294 7506
rect 25178 7394 25206 7506
rect 24266 7366 24670 7394
rect 24178 7254 24206 7366
rect 24642 7254 24670 7366
rect 24802 7366 25206 7394
rect 25250 7394 25278 7506
rect 25442 7394 25470 7506
rect 25250 7366 25294 7394
rect 24802 7254 24830 7366
rect 25266 7254 25294 7366
rect 25426 7366 25470 7394
rect 25514 7394 25542 7506
rect 26426 7394 26454 7506
rect 25514 7366 25918 7394
rect 25426 7254 25454 7366
rect 25890 7254 25918 7366
rect 26050 7366 26454 7394
rect 26498 7394 26526 7506
rect 26690 7394 26718 7506
rect 26498 7366 26542 7394
rect 26050 7254 26078 7366
rect 26514 7254 26542 7366
rect 26674 7366 26718 7394
rect 26762 7394 26790 7506
rect 27674 7394 27702 7506
rect 26762 7366 27166 7394
rect 26674 7254 26702 7366
rect 27138 7254 27166 7366
rect 27298 7366 27702 7394
rect 27746 7394 27774 7506
rect 27938 7394 27966 7506
rect 27746 7366 27790 7394
rect 27298 7254 27326 7366
rect 27762 7254 27790 7366
rect 27922 7366 27966 7394
rect 28010 7394 28038 7506
rect 28922 7394 28950 7506
rect 28010 7366 28414 7394
rect 27922 7254 27950 7366
rect 28386 7254 28414 7366
rect 28546 7366 28950 7394
rect 28994 7394 29022 7506
rect 29186 7394 29214 7506
rect 28994 7366 29038 7394
rect 28546 7254 28574 7366
rect 29010 7254 29038 7366
rect 29170 7366 29214 7394
rect 29258 7394 29286 7506
rect 30170 7394 30198 7506
rect 29258 7366 29662 7394
rect 29170 7254 29198 7366
rect 29634 7254 29662 7366
rect 29794 7366 30198 7394
rect 30242 7394 30270 7506
rect 30434 7394 30462 7506
rect 30242 7366 30286 7394
rect 29794 7254 29822 7366
rect 30258 7254 30286 7366
rect 30418 7366 30462 7394
rect 30506 7394 30534 7506
rect 31418 7394 31446 7506
rect 30506 7366 30910 7394
rect 30418 7254 30446 7366
rect 30882 7254 30910 7366
rect 31042 7366 31446 7394
rect 31490 7394 31518 7506
rect 31682 7394 31710 7506
rect 31490 7366 31534 7394
rect 31042 7254 31070 7366
rect 31506 7254 31534 7366
rect 31666 7366 31710 7394
rect 31754 7394 31782 7506
rect 32666 7394 32694 7506
rect 31754 7366 32158 7394
rect 31666 7254 31694 7366
rect 32130 7254 32158 7366
rect 32290 7366 32694 7394
rect 32738 7394 32766 7506
rect 32738 7366 32782 7394
rect 32290 7254 32318 7366
rect 32754 7254 32782 7366
rect 12786 6434 12814 6532
rect 12768 6382 12774 6434
rect 12826 6382 12832 6434
rect 6284 5043 6290 5095
rect 6342 5043 6348 5095
rect 6284 3553 6290 3605
rect 6342 3553 6348 3605
rect 4356 2212 4402 2270
rect 6284 2215 6290 2267
rect 6342 2215 6348 2267
rect 10571 1915 10577 1967
rect 10629 1955 10635 1967
rect 10629 1927 20907 1955
rect 10629 1915 10635 1927
rect 13103 1837 13163 1893
rect 15599 1837 15659 1893
rect 18095 1837 18155 1893
rect 20591 1837 20651 1893
rect 23087 1837 23147 1893
rect 25583 1837 25643 1893
rect 28079 1837 28139 1893
rect 30575 1837 30635 1893
rect 4232 722 4278 780
rect 6284 725 6290 777
rect 6342 725 6348 777
<< via1 >>
rect 39386 41188 39438 41197
rect 39386 41154 39395 41188
rect 39395 41154 39429 41188
rect 39429 41154 39438 41188
rect 39386 41145 39438 41154
rect 39386 39698 39438 39707
rect 39386 39664 39395 39698
rect 39395 39664 39429 39698
rect 39429 39664 39438 39698
rect 39386 39655 39438 39664
rect 39386 38360 39438 38369
rect 39386 38326 39395 38360
rect 39395 38326 39429 38360
rect 39429 38326 39438 38360
rect 39386 38317 39438 38326
rect 39386 36870 39438 36879
rect 39386 36836 39395 36870
rect 39395 36836 39429 36870
rect 39429 36836 39438 36870
rect 39386 36827 39438 36836
rect 32902 35488 32954 35540
rect 34868 33763 34920 33772
rect 34868 33729 34877 33763
rect 34877 33729 34911 33763
rect 34911 33729 34920 33763
rect 34868 33720 34920 33729
rect 10808 33523 10860 33532
rect 10808 33489 10817 33523
rect 10817 33489 10851 33523
rect 10851 33489 10860 33523
rect 10808 33480 10860 33489
rect 34868 33523 34920 33532
rect 34868 33489 34877 33523
rect 34877 33489 34911 33523
rect 34911 33489 34920 33523
rect 34868 33480 34920 33489
rect 10808 32973 10860 32982
rect 10808 32939 10817 32973
rect 10817 32939 10851 32973
rect 10851 32939 10860 32973
rect 10808 32930 10860 32939
rect 34868 32973 34920 32982
rect 34868 32939 34877 32973
rect 34877 32939 34911 32973
rect 34911 32939 34920 32973
rect 34868 32930 34920 32939
rect 10808 32733 10860 32742
rect 10808 32699 10817 32733
rect 10817 32699 10851 32733
rect 10851 32699 10860 32733
rect 10808 32690 10860 32699
rect 34868 32733 34920 32742
rect 34868 32699 34877 32733
rect 34877 32699 34911 32733
rect 34911 32699 34920 32733
rect 34868 32690 34920 32699
rect 10808 32183 10860 32192
rect 10808 32149 10817 32183
rect 10817 32149 10851 32183
rect 10851 32149 10860 32183
rect 10808 32140 10860 32149
rect 34868 32183 34920 32192
rect 34868 32149 34877 32183
rect 34877 32149 34911 32183
rect 34911 32149 34920 32183
rect 34868 32140 34920 32149
rect 10808 31943 10860 31952
rect 10808 31909 10817 31943
rect 10817 31909 10851 31943
rect 10851 31909 10860 31943
rect 10808 31900 10860 31909
rect 34868 31943 34920 31952
rect 34868 31909 34877 31943
rect 34877 31909 34911 31943
rect 34911 31909 34920 31943
rect 34868 31900 34920 31909
rect 10808 31393 10860 31402
rect 10808 31359 10817 31393
rect 10817 31359 10851 31393
rect 10851 31359 10860 31393
rect 10808 31350 10860 31359
rect 34868 31393 34920 31402
rect 34868 31359 34877 31393
rect 34877 31359 34911 31393
rect 34911 31359 34920 31393
rect 34868 31350 34920 31359
rect 10808 31153 10860 31162
rect 10808 31119 10817 31153
rect 10817 31119 10851 31153
rect 10851 31119 10860 31153
rect 10808 31110 10860 31119
rect 34868 31153 34920 31162
rect 34868 31119 34877 31153
rect 34877 31119 34911 31153
rect 34911 31119 34920 31153
rect 34868 31110 34920 31119
rect 10808 30603 10860 30612
rect 10808 30569 10817 30603
rect 10817 30569 10851 30603
rect 10851 30569 10860 30603
rect 10808 30560 10860 30569
rect 34868 30603 34920 30612
rect 34868 30569 34877 30603
rect 34877 30569 34911 30603
rect 34911 30569 34920 30603
rect 34868 30560 34920 30569
rect 10808 30363 10860 30372
rect 10808 30329 10817 30363
rect 10817 30329 10851 30363
rect 10851 30329 10860 30363
rect 10808 30320 10860 30329
rect 34868 30363 34920 30372
rect 34868 30329 34877 30363
rect 34877 30329 34911 30363
rect 34911 30329 34920 30363
rect 34868 30320 34920 30329
rect 10808 29813 10860 29822
rect 10808 29779 10817 29813
rect 10817 29779 10851 29813
rect 10851 29779 10860 29813
rect 10808 29770 10860 29779
rect 34868 29813 34920 29822
rect 34868 29779 34877 29813
rect 34877 29779 34911 29813
rect 34911 29779 34920 29813
rect 34868 29770 34920 29779
rect 10808 29573 10860 29582
rect 10808 29539 10817 29573
rect 10817 29539 10851 29573
rect 10851 29539 10860 29573
rect 10808 29530 10860 29539
rect 34868 29573 34920 29582
rect 34868 29539 34877 29573
rect 34877 29539 34911 29573
rect 34911 29539 34920 29573
rect 34868 29530 34920 29539
rect 10808 29023 10860 29032
rect 10808 28989 10817 29023
rect 10817 28989 10851 29023
rect 10851 28989 10860 29023
rect 10808 28980 10860 28989
rect 34868 29023 34920 29032
rect 34868 28989 34877 29023
rect 34877 28989 34911 29023
rect 34911 28989 34920 29023
rect 34868 28980 34920 28989
rect 10808 28783 10860 28792
rect 10808 28749 10817 28783
rect 10817 28749 10851 28783
rect 10851 28749 10860 28783
rect 10808 28740 10860 28749
rect 34868 28783 34920 28792
rect 34868 28749 34877 28783
rect 34877 28749 34911 28783
rect 34911 28749 34920 28783
rect 34868 28740 34920 28749
rect 10808 28233 10860 28242
rect 10808 28199 10817 28233
rect 10817 28199 10851 28233
rect 10851 28199 10860 28233
rect 10808 28190 10860 28199
rect 34868 28233 34920 28242
rect 34868 28199 34877 28233
rect 34877 28199 34911 28233
rect 34911 28199 34920 28233
rect 34868 28190 34920 28199
rect 10808 27993 10860 28002
rect 10808 27959 10817 27993
rect 10817 27959 10851 27993
rect 10851 27959 10860 27993
rect 10808 27950 10860 27959
rect 34868 27993 34920 28002
rect 34868 27959 34877 27993
rect 34877 27959 34911 27993
rect 34911 27959 34920 27993
rect 34868 27950 34920 27959
rect 10808 27443 10860 27452
rect 10808 27409 10817 27443
rect 10817 27409 10851 27443
rect 10851 27409 10860 27443
rect 10808 27400 10860 27409
rect 34868 27443 34920 27452
rect 34868 27409 34877 27443
rect 34877 27409 34911 27443
rect 34911 27409 34920 27443
rect 34868 27400 34920 27409
rect 10808 27203 10860 27212
rect 10808 27169 10817 27203
rect 10817 27169 10851 27203
rect 10851 27169 10860 27203
rect 10808 27160 10860 27169
rect 34868 27203 34920 27212
rect 34868 27169 34877 27203
rect 34877 27169 34911 27203
rect 34911 27169 34920 27203
rect 34868 27160 34920 27169
rect 10808 26653 10860 26662
rect 10808 26619 10817 26653
rect 10817 26619 10851 26653
rect 10851 26619 10860 26653
rect 10808 26610 10860 26619
rect 34868 26653 34920 26662
rect 34868 26619 34877 26653
rect 34877 26619 34911 26653
rect 34911 26619 34920 26653
rect 34868 26610 34920 26619
rect 10808 26413 10860 26422
rect 10808 26379 10817 26413
rect 10817 26379 10851 26413
rect 10851 26379 10860 26413
rect 10808 26370 10860 26379
rect 34868 26413 34920 26422
rect 34868 26379 34877 26413
rect 34877 26379 34911 26413
rect 34911 26379 34920 26413
rect 34868 26370 34920 26379
rect 10808 25863 10860 25872
rect 10808 25829 10817 25863
rect 10817 25829 10851 25863
rect 10851 25829 10860 25863
rect 10808 25820 10860 25829
rect 34868 25863 34920 25872
rect 34868 25829 34877 25863
rect 34877 25829 34911 25863
rect 34911 25829 34920 25863
rect 34868 25820 34920 25829
rect 10808 25623 10860 25632
rect 10808 25589 10817 25623
rect 10817 25589 10851 25623
rect 10851 25589 10860 25623
rect 10808 25580 10860 25589
rect 34868 25623 34920 25632
rect 34868 25589 34877 25623
rect 34877 25589 34911 25623
rect 34911 25589 34920 25623
rect 34868 25580 34920 25589
rect 10808 25073 10860 25082
rect 10808 25039 10817 25073
rect 10817 25039 10851 25073
rect 10851 25039 10860 25073
rect 10808 25030 10860 25039
rect 34868 25073 34920 25082
rect 34868 25039 34877 25073
rect 34877 25039 34911 25073
rect 34911 25039 34920 25073
rect 34868 25030 34920 25039
rect 10808 24833 10860 24842
rect 10808 24799 10817 24833
rect 10817 24799 10851 24833
rect 10851 24799 10860 24833
rect 10808 24790 10860 24799
rect 34868 24833 34920 24842
rect 34868 24799 34877 24833
rect 34877 24799 34911 24833
rect 34911 24799 34920 24833
rect 34868 24790 34920 24799
rect 10808 24283 10860 24292
rect 10808 24249 10817 24283
rect 10817 24249 10851 24283
rect 10851 24249 10860 24283
rect 10808 24240 10860 24249
rect 34868 24283 34920 24292
rect 34868 24249 34877 24283
rect 34877 24249 34911 24283
rect 34911 24249 34920 24283
rect 34868 24240 34920 24249
rect 10808 24043 10860 24052
rect 10808 24009 10817 24043
rect 10817 24009 10851 24043
rect 10851 24009 10860 24043
rect 10808 24000 10860 24009
rect 34868 24043 34920 24052
rect 34868 24009 34877 24043
rect 34877 24009 34911 24043
rect 34911 24009 34920 24043
rect 34868 24000 34920 24009
rect 10808 23493 10860 23502
rect 10808 23459 10817 23493
rect 10817 23459 10851 23493
rect 10851 23459 10860 23493
rect 10808 23450 10860 23459
rect 34868 23493 34920 23502
rect 34868 23459 34877 23493
rect 34877 23459 34911 23493
rect 34911 23459 34920 23493
rect 34868 23450 34920 23459
rect 10808 23253 10860 23262
rect 10808 23219 10817 23253
rect 10817 23219 10851 23253
rect 10851 23219 10860 23253
rect 10808 23210 10860 23219
rect 34868 23253 34920 23262
rect 34868 23219 34877 23253
rect 34877 23219 34911 23253
rect 34911 23219 34920 23253
rect 34868 23210 34920 23219
rect 10808 22703 10860 22712
rect 10808 22669 10817 22703
rect 10817 22669 10851 22703
rect 10851 22669 10860 22703
rect 10808 22660 10860 22669
rect 34868 22703 34920 22712
rect 34868 22669 34877 22703
rect 34877 22669 34911 22703
rect 34911 22669 34920 22703
rect 34868 22660 34920 22669
rect 10808 22463 10860 22472
rect 10808 22429 10817 22463
rect 10817 22429 10851 22463
rect 10851 22429 10860 22463
rect 10808 22420 10860 22429
rect 34868 22463 34920 22472
rect 34868 22429 34877 22463
rect 34877 22429 34911 22463
rect 34911 22429 34920 22463
rect 34868 22420 34920 22429
rect 10808 21913 10860 21922
rect 10808 21879 10817 21913
rect 10817 21879 10851 21913
rect 10851 21879 10860 21913
rect 10808 21870 10860 21879
rect 34868 21913 34920 21922
rect 34868 21879 34877 21913
rect 34877 21879 34911 21913
rect 34911 21879 34920 21913
rect 34868 21870 34920 21879
rect 10808 21673 10860 21682
rect 10808 21639 10817 21673
rect 10817 21639 10851 21673
rect 10851 21639 10860 21673
rect 10808 21630 10860 21639
rect 34868 21673 34920 21682
rect 34868 21639 34877 21673
rect 34877 21639 34911 21673
rect 34911 21639 34920 21673
rect 34868 21630 34920 21639
rect 10808 21123 10860 21132
rect 10808 21089 10817 21123
rect 10817 21089 10851 21123
rect 10851 21089 10860 21123
rect 10808 21080 10860 21089
rect 34868 21123 34920 21132
rect 34868 21089 34877 21123
rect 34877 21089 34911 21123
rect 34911 21089 34920 21123
rect 34868 21080 34920 21089
rect 10808 20883 10860 20892
rect 10808 20849 10817 20883
rect 10817 20849 10851 20883
rect 10851 20849 10860 20883
rect 10808 20840 10860 20849
rect 34868 20883 34920 20892
rect 34868 20849 34877 20883
rect 34877 20849 34911 20883
rect 34911 20849 34920 20883
rect 34868 20840 34920 20849
rect 10808 20333 10860 20342
rect 10808 20299 10817 20333
rect 10817 20299 10851 20333
rect 10851 20299 10860 20333
rect 10808 20290 10860 20299
rect 34868 20333 34920 20342
rect 34868 20299 34877 20333
rect 34877 20299 34911 20333
rect 34911 20299 34920 20333
rect 34868 20290 34920 20299
rect 10808 20093 10860 20102
rect 10808 20059 10817 20093
rect 10817 20059 10851 20093
rect 10851 20059 10860 20093
rect 10808 20050 10860 20059
rect 34868 20093 34920 20102
rect 34868 20059 34877 20093
rect 34877 20059 34911 20093
rect 34911 20059 34920 20093
rect 34868 20050 34920 20059
rect 10808 19543 10860 19552
rect 10808 19509 10817 19543
rect 10817 19509 10851 19543
rect 10851 19509 10860 19543
rect 10808 19500 10860 19509
rect 34868 19543 34920 19552
rect 34868 19509 34877 19543
rect 34877 19509 34911 19543
rect 34911 19509 34920 19543
rect 34868 19500 34920 19509
rect 10808 19303 10860 19312
rect 10808 19269 10817 19303
rect 10817 19269 10851 19303
rect 10851 19269 10860 19303
rect 10808 19260 10860 19269
rect 34868 19303 34920 19312
rect 34868 19269 34877 19303
rect 34877 19269 34911 19303
rect 34911 19269 34920 19303
rect 34868 19260 34920 19269
rect 10808 18753 10860 18762
rect 10808 18719 10817 18753
rect 10817 18719 10851 18753
rect 10851 18719 10860 18753
rect 10808 18710 10860 18719
rect 34868 18753 34920 18762
rect 34868 18719 34877 18753
rect 34877 18719 34911 18753
rect 34911 18719 34920 18753
rect 34868 18710 34920 18719
rect 10808 18513 10860 18522
rect 10808 18479 10817 18513
rect 10817 18479 10851 18513
rect 10851 18479 10860 18513
rect 10808 18470 10860 18479
rect 34868 18513 34920 18522
rect 34868 18479 34877 18513
rect 34877 18479 34911 18513
rect 34911 18479 34920 18513
rect 34868 18470 34920 18479
rect 10808 17963 10860 17972
rect 10808 17929 10817 17963
rect 10817 17929 10851 17963
rect 10851 17929 10860 17963
rect 10808 17920 10860 17929
rect 34868 17963 34920 17972
rect 34868 17929 34877 17963
rect 34877 17929 34911 17963
rect 34911 17929 34920 17963
rect 34868 17920 34920 17929
rect 10808 17723 10860 17732
rect 10808 17689 10817 17723
rect 10817 17689 10851 17723
rect 10851 17689 10860 17723
rect 10808 17680 10860 17689
rect 34868 17723 34920 17732
rect 34868 17689 34877 17723
rect 34877 17689 34911 17723
rect 34911 17689 34920 17723
rect 34868 17680 34920 17689
rect 10808 17173 10860 17182
rect 10808 17139 10817 17173
rect 10817 17139 10851 17173
rect 10851 17139 10860 17173
rect 10808 17130 10860 17139
rect 34868 17173 34920 17182
rect 34868 17139 34877 17173
rect 34877 17139 34911 17173
rect 34911 17139 34920 17173
rect 34868 17130 34920 17139
rect 10808 16933 10860 16942
rect 10808 16899 10817 16933
rect 10817 16899 10851 16933
rect 10851 16899 10860 16933
rect 10808 16890 10860 16899
rect 34868 16933 34920 16942
rect 34868 16899 34877 16933
rect 34877 16899 34911 16933
rect 34911 16899 34920 16933
rect 34868 16890 34920 16899
rect 10808 16383 10860 16392
rect 10808 16349 10817 16383
rect 10817 16349 10851 16383
rect 10851 16349 10860 16383
rect 10808 16340 10860 16349
rect 34868 16383 34920 16392
rect 34868 16349 34877 16383
rect 34877 16349 34911 16383
rect 34911 16349 34920 16383
rect 34868 16340 34920 16349
rect 10808 16143 10860 16152
rect 10808 16109 10817 16143
rect 10817 16109 10851 16143
rect 10851 16109 10860 16143
rect 10808 16100 10860 16109
rect 34868 16143 34920 16152
rect 34868 16109 34877 16143
rect 34877 16109 34911 16143
rect 34911 16109 34920 16143
rect 34868 16100 34920 16109
rect 10808 15593 10860 15602
rect 10808 15559 10817 15593
rect 10817 15559 10851 15593
rect 10851 15559 10860 15593
rect 10808 15550 10860 15559
rect 34868 15593 34920 15602
rect 34868 15559 34877 15593
rect 34877 15559 34911 15593
rect 34911 15559 34920 15593
rect 34868 15550 34920 15559
rect 10808 15353 10860 15362
rect 10808 15319 10817 15353
rect 10817 15319 10851 15353
rect 10851 15319 10860 15353
rect 10808 15310 10860 15319
rect 34868 15353 34920 15362
rect 34868 15319 34877 15353
rect 34877 15319 34911 15353
rect 34911 15319 34920 15353
rect 34868 15310 34920 15319
rect 10808 14803 10860 14812
rect 10808 14769 10817 14803
rect 10817 14769 10851 14803
rect 10851 14769 10860 14803
rect 10808 14760 10860 14769
rect 34868 14803 34920 14812
rect 34868 14769 34877 14803
rect 34877 14769 34911 14803
rect 34911 14769 34920 14803
rect 34868 14760 34920 14769
rect 10808 14563 10860 14572
rect 10808 14529 10817 14563
rect 10817 14529 10851 14563
rect 10851 14529 10860 14563
rect 10808 14520 10860 14529
rect 34868 14563 34920 14572
rect 34868 14529 34877 14563
rect 34877 14529 34911 14563
rect 34911 14529 34920 14563
rect 34868 14520 34920 14529
rect 10808 14013 10860 14022
rect 10808 13979 10817 14013
rect 10817 13979 10851 14013
rect 10851 13979 10860 14013
rect 10808 13970 10860 13979
rect 34868 14013 34920 14022
rect 34868 13979 34877 14013
rect 34877 13979 34911 14013
rect 34911 13979 34920 14013
rect 34868 13970 34920 13979
rect 10808 13773 10860 13782
rect 10808 13739 10817 13773
rect 10817 13739 10851 13773
rect 10851 13739 10860 13773
rect 10808 13730 10860 13739
rect 34868 13773 34920 13782
rect 34868 13739 34877 13773
rect 34877 13739 34911 13773
rect 34911 13739 34920 13773
rect 34868 13730 34920 13739
rect 10808 13223 10860 13232
rect 10808 13189 10817 13223
rect 10817 13189 10851 13223
rect 10851 13189 10860 13223
rect 10808 13180 10860 13189
rect 34868 13223 34920 13232
rect 34868 13189 34877 13223
rect 34877 13189 34911 13223
rect 34911 13189 34920 13223
rect 34868 13180 34920 13189
rect 10808 12983 10860 12992
rect 10808 12949 10817 12983
rect 10817 12949 10851 12983
rect 10851 12949 10860 12983
rect 10808 12940 10860 12949
rect 34868 12983 34920 12992
rect 34868 12949 34877 12983
rect 34877 12949 34911 12983
rect 34911 12949 34920 12983
rect 34868 12940 34920 12949
rect 10808 12433 10860 12442
rect 10808 12399 10817 12433
rect 10817 12399 10851 12433
rect 10851 12399 10860 12433
rect 10808 12390 10860 12399
rect 34868 12433 34920 12442
rect 34868 12399 34877 12433
rect 34877 12399 34911 12433
rect 34911 12399 34920 12433
rect 34868 12390 34920 12399
rect 10808 12193 10860 12202
rect 10808 12159 10817 12193
rect 10817 12159 10851 12193
rect 10851 12159 10860 12193
rect 10808 12150 10860 12159
rect 34868 12193 34920 12202
rect 34868 12159 34877 12193
rect 34877 12159 34911 12193
rect 34911 12159 34920 12193
rect 34868 12150 34920 12159
rect 10808 11643 10860 11652
rect 10808 11609 10817 11643
rect 10817 11609 10851 11643
rect 10851 11609 10860 11643
rect 10808 11600 10860 11609
rect 34868 11643 34920 11652
rect 34868 11609 34877 11643
rect 34877 11609 34911 11643
rect 34911 11609 34920 11643
rect 34868 11600 34920 11609
rect 10808 11403 10860 11412
rect 10808 11369 10817 11403
rect 10817 11369 10851 11403
rect 10851 11369 10860 11403
rect 10808 11360 10860 11369
rect 34868 11403 34920 11412
rect 34868 11369 34877 11403
rect 34877 11369 34911 11403
rect 34911 11369 34920 11403
rect 34868 11360 34920 11369
rect 10808 10853 10860 10862
rect 10808 10819 10817 10853
rect 10817 10819 10851 10853
rect 10851 10819 10860 10853
rect 10808 10810 10860 10819
rect 34868 10853 34920 10862
rect 34868 10819 34877 10853
rect 34877 10819 34911 10853
rect 34911 10819 34920 10853
rect 34868 10810 34920 10819
rect 10808 10613 10860 10622
rect 10808 10579 10817 10613
rect 10817 10579 10851 10613
rect 10851 10579 10860 10613
rect 10808 10570 10860 10579
rect 34868 10613 34920 10622
rect 34868 10579 34877 10613
rect 34877 10579 34911 10613
rect 34911 10579 34920 10613
rect 34868 10570 34920 10579
rect 10808 10063 10860 10072
rect 10808 10029 10817 10063
rect 10817 10029 10851 10063
rect 10851 10029 10860 10063
rect 10808 10020 10860 10029
rect 34868 10063 34920 10072
rect 34868 10029 34877 10063
rect 34877 10029 34911 10063
rect 34911 10029 34920 10063
rect 34868 10020 34920 10029
rect 10808 9823 10860 9832
rect 10808 9789 10817 9823
rect 10817 9789 10851 9823
rect 10851 9789 10860 9823
rect 10808 9780 10860 9789
rect 34868 9823 34920 9832
rect 34868 9789 34877 9823
rect 34877 9789 34911 9823
rect 34911 9789 34920 9823
rect 34868 9780 34920 9789
rect 10808 9273 10860 9282
rect 10808 9239 10817 9273
rect 10817 9239 10851 9273
rect 10851 9239 10860 9273
rect 10808 9230 10860 9239
rect 34868 9273 34920 9282
rect 34868 9239 34877 9273
rect 34877 9239 34911 9273
rect 34911 9239 34920 9273
rect 34868 9230 34920 9239
rect 10808 9033 10860 9042
rect 10808 8999 10817 9033
rect 10817 8999 10851 9033
rect 10851 8999 10860 9033
rect 10808 8990 10860 8999
rect 34868 9033 34920 9042
rect 34868 8999 34877 9033
rect 34877 8999 34911 9033
rect 34911 8999 34920 9033
rect 34868 8990 34920 8999
rect 10808 8483 10860 8492
rect 10808 8449 10817 8483
rect 10817 8449 10851 8483
rect 10851 8449 10860 8483
rect 10808 8440 10860 8449
rect 34868 8483 34920 8492
rect 34868 8449 34877 8483
rect 34877 8449 34911 8483
rect 34911 8449 34920 8483
rect 34868 8440 34920 8449
rect 10808 8243 10860 8252
rect 10808 8209 10817 8243
rect 10817 8209 10851 8243
rect 10851 8209 10860 8243
rect 10808 8200 10860 8209
rect 12774 6382 12826 6434
rect 6290 5086 6342 5095
rect 6290 5052 6299 5086
rect 6299 5052 6333 5086
rect 6333 5052 6342 5086
rect 6290 5043 6342 5052
rect 6290 3596 6342 3605
rect 6290 3562 6299 3596
rect 6299 3562 6333 3596
rect 6333 3562 6342 3596
rect 6290 3553 6342 3562
rect 6290 2258 6342 2267
rect 6290 2224 6299 2258
rect 6299 2224 6333 2258
rect 6333 2224 6342 2258
rect 6290 2215 6342 2224
rect 10577 1915 10629 1967
rect 6290 768 6342 777
rect 6290 734 6299 768
rect 6299 734 6333 768
rect 6333 734 6342 768
rect 6290 725 6342 734
<< metal2 >>
rect 35077 38177 35105 41924
rect 35063 38168 35119 38177
rect 35063 38103 35119 38112
rect 32900 35542 32956 35551
rect 32900 35477 32956 35486
rect 35077 34416 35105 38103
rect 35201 35402 35229 41924
rect 38881 41199 38937 41208
rect 38881 41134 38937 41143
rect 39384 41199 39440 41208
rect 39384 41134 39440 41143
rect 38609 39709 38665 39718
rect 38609 39644 38665 39653
rect 38623 37337 38651 39644
rect 38745 38371 38801 38380
rect 38745 38306 38801 38315
rect 38609 37328 38665 37337
rect 38609 37263 38665 37272
rect 38759 37213 38787 38306
rect 38895 37461 38923 41134
rect 39384 39709 39440 39718
rect 39384 39644 39440 39653
rect 39384 38371 39440 38380
rect 39384 38306 39440 38315
rect 38881 37452 38937 37461
rect 38881 37387 38937 37396
rect 38745 37204 38801 37213
rect 38745 37139 38801 37148
rect 38609 37080 38665 37089
rect 38609 37015 38665 37024
rect 38623 36890 38651 37015
rect 38609 36881 38665 36890
rect 38609 36816 38665 36825
rect 39384 36881 39440 36890
rect 39384 36816 39440 36825
rect 35187 35393 35243 35402
rect 35187 35328 35243 35337
rect 35201 34416 35229 35328
rect 38262 33911 38290 33939
rect 34868 33772 34920 33778
rect 34146 33739 34868 33767
rect 34868 33714 34920 33720
rect 10808 33532 10860 33538
rect 34868 33532 34920 33538
rect 34146 33485 34868 33513
rect 10808 33474 10860 33480
rect 34868 33474 34920 33480
rect 10820 33293 10848 33474
rect 10820 33265 11582 33293
rect 10820 33169 11582 33197
rect 10820 32988 10848 33169
rect 10808 32982 10860 32988
rect 34868 32982 34920 32988
rect 34146 32949 34868 32977
rect 10808 32924 10860 32930
rect 34868 32924 34920 32930
rect 10808 32742 10860 32748
rect 34868 32742 34920 32748
rect 34146 32695 34868 32723
rect 10808 32684 10860 32690
rect 34868 32684 34920 32690
rect 10820 32503 10848 32684
rect 10820 32475 11582 32503
rect 10820 32379 11582 32407
rect 10820 32198 10848 32379
rect 10808 32192 10860 32198
rect 34868 32192 34920 32198
rect 34146 32159 34868 32187
rect 10808 32134 10860 32140
rect 34868 32134 34920 32140
rect 10808 31952 10860 31958
rect 34868 31952 34920 31958
rect 34146 31905 34868 31933
rect 10808 31894 10860 31900
rect 34868 31894 34920 31900
rect 10820 31713 10848 31894
rect 10820 31685 11582 31713
rect 10820 31589 11582 31617
rect 10820 31408 10848 31589
rect 10808 31402 10860 31408
rect 34868 31402 34920 31408
rect 34146 31369 34868 31397
rect 10808 31344 10860 31350
rect 34868 31344 34920 31350
rect 10808 31162 10860 31168
rect 34868 31162 34920 31168
rect 34146 31115 34868 31143
rect 10808 31104 10860 31110
rect 34868 31104 34920 31110
rect 10820 30923 10848 31104
rect 10820 30895 11582 30923
rect 10820 30799 11582 30827
rect 10820 30618 10848 30799
rect 10808 30612 10860 30618
rect 34868 30612 34920 30618
rect 34146 30579 34868 30607
rect 10808 30554 10860 30560
rect 34868 30554 34920 30560
rect 10808 30372 10860 30378
rect 34868 30372 34920 30378
rect 34146 30325 34868 30353
rect 10808 30314 10860 30320
rect 34868 30314 34920 30320
rect 10820 30133 10848 30314
rect 10820 30105 11582 30133
rect 10820 30009 11582 30037
rect 10820 29828 10848 30009
rect 10808 29822 10860 29828
rect 34868 29822 34920 29828
rect 34146 29789 34868 29817
rect 10808 29764 10860 29770
rect 34868 29764 34920 29770
rect 10808 29582 10860 29588
rect 34868 29582 34920 29588
rect 34146 29535 34868 29563
rect 10808 29524 10860 29530
rect 34868 29524 34920 29530
rect 10820 29343 10848 29524
rect 10820 29315 11582 29343
rect 10820 29219 11582 29247
rect 10820 29038 10848 29219
rect 10808 29032 10860 29038
rect 34868 29032 34920 29038
rect 34146 28999 34868 29027
rect 10808 28974 10860 28980
rect 34868 28974 34920 28980
rect 10808 28792 10860 28798
rect 34868 28792 34920 28798
rect 34146 28745 34868 28773
rect 10808 28734 10860 28740
rect 34868 28734 34920 28740
rect 10820 28553 10848 28734
rect 10820 28525 11582 28553
rect 10820 28429 11582 28457
rect 10820 28248 10848 28429
rect 10808 28242 10860 28248
rect 34868 28242 34920 28248
rect 34146 28209 34868 28237
rect 10808 28184 10860 28190
rect 34868 28184 34920 28190
rect 10808 28002 10860 28008
rect 34868 28002 34920 28008
rect 34146 27955 34868 27983
rect 10808 27944 10860 27950
rect 34868 27944 34920 27950
rect 10820 27763 10848 27944
rect 10820 27735 11582 27763
rect 10820 27639 11582 27667
rect 10820 27458 10848 27639
rect 10808 27452 10860 27458
rect 34868 27452 34920 27458
rect 34146 27419 34868 27447
rect 10808 27394 10860 27400
rect 34868 27394 34920 27400
rect 10808 27212 10860 27218
rect 34868 27212 34920 27218
rect 34146 27165 34868 27193
rect 10808 27154 10860 27160
rect 34868 27154 34920 27160
rect 10820 26973 10848 27154
rect 10820 26945 11582 26973
rect 10820 26849 11582 26877
rect 10820 26668 10848 26849
rect 10808 26662 10860 26668
rect 34868 26662 34920 26668
rect 34146 26629 34868 26657
rect 10808 26604 10860 26610
rect 34868 26604 34920 26610
rect 10808 26422 10860 26428
rect 34868 26422 34920 26428
rect 34146 26375 34868 26403
rect 10808 26364 10860 26370
rect 34868 26364 34920 26370
rect 10820 26183 10848 26364
rect 10820 26155 11582 26183
rect 10820 26059 11582 26087
rect 10820 25878 10848 26059
rect 10808 25872 10860 25878
rect 34868 25872 34920 25878
rect 34146 25839 34868 25867
rect 10808 25814 10860 25820
rect 34868 25814 34920 25820
rect 10808 25632 10860 25638
rect 34868 25632 34920 25638
rect 34146 25585 34868 25613
rect 10808 25574 10860 25580
rect 34868 25574 34920 25580
rect 10820 25393 10848 25574
rect 10820 25365 11582 25393
rect 10820 25269 11582 25297
rect 10820 25088 10848 25269
rect 10808 25082 10860 25088
rect 34868 25082 34920 25088
rect 34146 25049 34868 25077
rect 10808 25024 10860 25030
rect 34868 25024 34920 25030
rect 10808 24842 10860 24848
rect 34868 24842 34920 24848
rect 34146 24795 34868 24823
rect 10808 24784 10860 24790
rect 34868 24784 34920 24790
rect 10820 24603 10848 24784
rect 10820 24575 11582 24603
rect 10820 24479 11582 24507
rect 10820 24298 10848 24479
rect 10808 24292 10860 24298
rect 34868 24292 34920 24298
rect 34146 24259 34868 24287
rect 10808 24234 10860 24240
rect 34868 24234 34920 24240
rect 10808 24052 10860 24058
rect 34868 24052 34920 24058
rect 34146 24005 34868 24033
rect 10808 23994 10860 24000
rect 34868 23994 34920 24000
rect 10820 23813 10848 23994
rect 10820 23785 11582 23813
rect 10820 23689 11582 23717
rect 10820 23508 10848 23689
rect 10808 23502 10860 23508
rect 34868 23502 34920 23508
rect 34146 23469 34868 23497
rect 10808 23444 10860 23450
rect 34868 23444 34920 23450
rect 10808 23262 10860 23268
rect 34868 23262 34920 23268
rect 34146 23215 34868 23243
rect 10808 23204 10860 23210
rect 34868 23204 34920 23210
rect 10820 23023 10848 23204
rect 10820 22995 11582 23023
rect 10820 22899 11582 22927
rect 10820 22718 10848 22899
rect 10808 22712 10860 22718
rect 34868 22712 34920 22718
rect 34146 22679 34868 22707
rect 10808 22654 10860 22660
rect 34868 22654 34920 22660
rect 10808 22472 10860 22478
rect 34868 22472 34920 22478
rect 34146 22425 34868 22453
rect 10808 22414 10860 22420
rect 34868 22414 34920 22420
rect 10820 22233 10848 22414
rect 10820 22205 11582 22233
rect 10820 22109 11582 22137
rect 10820 21928 10848 22109
rect 10808 21922 10860 21928
rect 34868 21922 34920 21928
rect 34146 21889 34868 21917
rect 10808 21864 10860 21870
rect 34868 21864 34920 21870
rect 10808 21682 10860 21688
rect 34868 21682 34920 21688
rect 34146 21635 34868 21663
rect 10808 21624 10860 21630
rect 34868 21624 34920 21630
rect 10820 21443 10848 21624
rect 10820 21415 11582 21443
rect 10820 21319 11582 21347
rect 10820 21138 10848 21319
rect 10808 21132 10860 21138
rect 34868 21132 34920 21138
rect 34146 21099 34868 21127
rect 10808 21074 10860 21080
rect 34868 21074 34920 21080
rect 10808 20892 10860 20898
rect 34868 20892 34920 20898
rect 34146 20845 34868 20873
rect 10808 20834 10860 20840
rect 34868 20834 34920 20840
rect 10820 20653 10848 20834
rect 10820 20625 11582 20653
rect 10820 20529 11582 20557
rect 10820 20348 10848 20529
rect 10808 20342 10860 20348
rect 34868 20342 34920 20348
rect 34146 20309 34868 20337
rect 10808 20284 10860 20290
rect 34868 20284 34920 20290
rect 10808 20102 10860 20108
rect 34868 20102 34920 20108
rect 34146 20055 34868 20083
rect 10808 20044 10860 20050
rect 34868 20044 34920 20050
rect 10820 19863 10848 20044
rect 10820 19835 11582 19863
rect 10820 19739 11582 19767
rect 10820 19558 10848 19739
rect 10808 19552 10860 19558
rect 34868 19552 34920 19558
rect 34146 19519 34868 19547
rect 10808 19494 10860 19500
rect 34868 19494 34920 19500
rect 10808 19312 10860 19318
rect 34868 19312 34920 19318
rect 34146 19265 34868 19293
rect 10808 19254 10860 19260
rect 34868 19254 34920 19260
rect 10820 19073 10848 19254
rect 10820 19045 11582 19073
rect 10820 18949 11582 18977
rect 10820 18768 10848 18949
rect 10808 18762 10860 18768
rect 34868 18762 34920 18768
rect 34146 18729 34868 18757
rect 10808 18704 10860 18710
rect 34868 18704 34920 18710
rect 10808 18522 10860 18528
rect 34868 18522 34920 18528
rect 34146 18475 34868 18503
rect 10808 18464 10860 18470
rect 34868 18464 34920 18470
rect 10820 18283 10848 18464
rect 10820 18255 11582 18283
rect 10820 18159 11582 18187
rect 10820 17978 10848 18159
rect 10808 17972 10860 17978
rect 34868 17972 34920 17978
rect 34146 17939 34868 17967
rect 10808 17914 10860 17920
rect 34868 17914 34920 17920
rect 10808 17732 10860 17738
rect 34868 17732 34920 17738
rect 34146 17685 34868 17713
rect 10808 17674 10860 17680
rect 34868 17674 34920 17680
rect 10820 17493 10848 17674
rect 10820 17465 11582 17493
rect 10820 17369 11582 17397
rect 10820 17188 10848 17369
rect 10808 17182 10860 17188
rect 34868 17182 34920 17188
rect 34146 17149 34868 17177
rect 10808 17124 10860 17130
rect 34868 17124 34920 17130
rect 10808 16942 10860 16948
rect 34868 16942 34920 16948
rect 34146 16895 34868 16923
rect 10808 16884 10860 16890
rect 34868 16884 34920 16890
rect 10820 16703 10848 16884
rect 10820 16675 11582 16703
rect 10820 16579 11582 16607
rect 10820 16398 10848 16579
rect 10808 16392 10860 16398
rect 34868 16392 34920 16398
rect 34146 16359 34868 16387
rect 10808 16334 10860 16340
rect 34868 16334 34920 16340
rect 10808 16152 10860 16158
rect 34868 16152 34920 16158
rect 34146 16105 34868 16133
rect 10808 16094 10860 16100
rect 34868 16094 34920 16100
rect 10820 15913 10848 16094
rect 10820 15885 11582 15913
rect 10820 15789 11582 15817
rect 10820 15608 10848 15789
rect 10808 15602 10860 15608
rect 34868 15602 34920 15608
rect 34146 15569 34868 15597
rect 10808 15544 10860 15550
rect 34868 15544 34920 15550
rect 10808 15362 10860 15368
rect 34868 15362 34920 15368
rect 34146 15315 34868 15343
rect 10808 15304 10860 15310
rect 34868 15304 34920 15310
rect 10820 15123 10848 15304
rect 10820 15095 11582 15123
rect 10820 14999 11582 15027
rect 10820 14818 10848 14999
rect 10808 14812 10860 14818
rect 34868 14812 34920 14818
rect 34146 14779 34868 14807
rect 10808 14754 10860 14760
rect 34868 14754 34920 14760
rect 10808 14572 10860 14578
rect 34868 14572 34920 14578
rect 34146 14525 34868 14553
rect 10808 14514 10860 14520
rect 34868 14514 34920 14520
rect 10820 14333 10848 14514
rect 10820 14305 11582 14333
rect 10820 14209 11582 14237
rect 10820 14028 10848 14209
rect 10808 14022 10860 14028
rect 34868 14022 34920 14028
rect 34146 13989 34868 14017
rect 10808 13964 10860 13970
rect 34868 13964 34920 13970
rect 10808 13782 10860 13788
rect 34868 13782 34920 13788
rect 34146 13735 34868 13763
rect 10808 13724 10860 13730
rect 34868 13724 34920 13730
rect 10820 13543 10848 13724
rect 10820 13515 11582 13543
rect 10820 13419 11582 13447
rect 10820 13238 10848 13419
rect 10808 13232 10860 13238
rect 34868 13232 34920 13238
rect 34146 13199 34868 13227
rect 10808 13174 10860 13180
rect 34868 13174 34920 13180
rect 10808 12992 10860 12998
rect 34868 12992 34920 12998
rect 34146 12945 34868 12973
rect 10808 12934 10860 12940
rect 34868 12934 34920 12940
rect 10820 12753 10848 12934
rect 10820 12725 11582 12753
rect 10820 12629 11582 12657
rect 10820 12448 10848 12629
rect 10808 12442 10860 12448
rect 34868 12442 34920 12448
rect 34146 12409 34868 12437
rect 10808 12384 10860 12390
rect 34868 12384 34920 12390
rect 10808 12202 10860 12208
rect 34868 12202 34920 12208
rect 34146 12155 34868 12183
rect 10808 12144 10860 12150
rect 34868 12144 34920 12150
rect 10820 11963 10848 12144
rect 10820 11935 11582 11963
rect 10820 11839 11582 11867
rect 10820 11658 10848 11839
rect 10808 11652 10860 11658
rect 34868 11652 34920 11658
rect 34146 11619 34868 11647
rect 10808 11594 10860 11600
rect 34868 11594 34920 11600
rect 10808 11412 10860 11418
rect 34868 11412 34920 11418
rect 34146 11365 34868 11393
rect 10808 11354 10860 11360
rect 34868 11354 34920 11360
rect 10820 11173 10848 11354
rect 10820 11145 11582 11173
rect 10820 11049 11582 11077
rect 10820 10868 10848 11049
rect 10808 10862 10860 10868
rect 34868 10862 34920 10868
rect 34146 10829 34868 10857
rect 10808 10804 10860 10810
rect 34868 10804 34920 10810
rect 10808 10622 10860 10628
rect 34868 10622 34920 10628
rect 34146 10575 34868 10603
rect 10808 10564 10860 10570
rect 34868 10564 34920 10570
rect 10820 10383 10848 10564
rect 10820 10355 11582 10383
rect 10820 10259 11582 10287
rect 10820 10078 10848 10259
rect 10808 10072 10860 10078
rect 34868 10072 34920 10078
rect 34146 10039 34868 10067
rect 10808 10014 10860 10020
rect 34868 10014 34920 10020
rect 10808 9832 10860 9838
rect 34868 9832 34920 9838
rect 34146 9785 34868 9813
rect 10808 9774 10860 9780
rect 34868 9774 34920 9780
rect 10820 9593 10848 9774
rect 10820 9565 11582 9593
rect 10820 9469 11582 9497
rect 10820 9288 10848 9469
rect 10808 9282 10860 9288
rect 34868 9282 34920 9288
rect 34146 9249 34868 9277
rect 10808 9224 10860 9230
rect 34868 9224 34920 9230
rect 10808 9042 10860 9048
rect 34868 9042 34920 9048
rect 34146 8995 34868 9023
rect 10808 8984 10860 8990
rect 34868 8984 34920 8990
rect 10820 8803 10848 8984
rect 10820 8775 11582 8803
rect 10820 8679 11582 8707
rect 10820 8498 10848 8679
rect 10808 8492 10860 8498
rect 34868 8492 34920 8498
rect 34146 8459 34868 8487
rect 10808 8434 10860 8440
rect 34868 8434 34920 8440
rect 10808 8252 10860 8258
rect 10808 8194 10860 8200
rect 7438 8033 7466 8061
rect 10820 8013 10848 8194
rect 10820 7985 11582 8013
rect 10465 6594 10493 7506
rect 10451 6585 10507 6594
rect 10451 6520 10507 6529
rect 6288 5097 6344 5106
rect 6288 5032 6344 5041
rect 6567 5097 6623 5106
rect 6567 5032 6623 5041
rect 6581 4907 6609 5032
rect 6567 4898 6623 4907
rect 6567 4833 6623 4842
rect 6839 4774 6895 4783
rect 6839 4709 6895 4718
rect 6703 4650 6759 4659
rect 6703 4585 6759 4594
rect 6567 4526 6623 4535
rect 6567 4461 6623 4470
rect 6288 3607 6344 3616
rect 6288 3542 6344 3551
rect 6288 2269 6344 2278
rect 6288 2204 6344 2213
rect 6581 788 6609 4461
rect 6717 2278 6745 4585
rect 6853 3616 6881 4709
rect 6839 3607 6895 3616
rect 6839 3542 6895 3551
rect 6703 2269 6759 2278
rect 6703 2204 6759 2213
rect 6288 779 6344 788
rect 6288 714 6344 723
rect 6567 779 6623 788
rect 6567 714 6623 723
rect 10465 82 10493 6520
rect 10589 1973 10617 7506
rect 12772 6436 12828 6445
rect 12772 6371 12828 6380
rect 10577 1967 10629 1973
rect 10577 1909 10629 1915
rect 10589 82 10617 1909
<< via2 >>
rect 35063 38112 35119 38168
rect 32900 35540 32956 35542
rect 32900 35488 32902 35540
rect 32902 35488 32954 35540
rect 32954 35488 32956 35540
rect 32900 35486 32956 35488
rect 38881 41143 38937 41199
rect 39384 41197 39440 41199
rect 39384 41145 39386 41197
rect 39386 41145 39438 41197
rect 39438 41145 39440 41197
rect 39384 41143 39440 41145
rect 38609 39653 38665 39709
rect 38745 38315 38801 38371
rect 38609 37272 38665 37328
rect 39384 39707 39440 39709
rect 39384 39655 39386 39707
rect 39386 39655 39438 39707
rect 39438 39655 39440 39707
rect 39384 39653 39440 39655
rect 39384 38369 39440 38371
rect 39384 38317 39386 38369
rect 39386 38317 39438 38369
rect 39438 38317 39440 38369
rect 39384 38315 39440 38317
rect 38881 37396 38937 37452
rect 38745 37148 38801 37204
rect 38609 37024 38665 37080
rect 38609 36825 38665 36881
rect 39384 36879 39440 36881
rect 39384 36827 39386 36879
rect 39386 36827 39438 36879
rect 39438 36827 39440 36879
rect 39384 36825 39440 36827
rect 35187 35337 35243 35393
rect 10451 6529 10507 6585
rect 6288 5095 6344 5097
rect 6288 5043 6290 5095
rect 6290 5043 6342 5095
rect 6342 5043 6344 5095
rect 6288 5041 6344 5043
rect 6567 5041 6623 5097
rect 6567 4842 6623 4898
rect 6839 4718 6895 4774
rect 6703 4594 6759 4650
rect 6567 4470 6623 4526
rect 6288 3605 6344 3607
rect 6288 3553 6290 3605
rect 6290 3553 6342 3605
rect 6342 3553 6344 3605
rect 6288 3551 6344 3553
rect 6288 2267 6344 2269
rect 6288 2215 6290 2267
rect 6290 2215 6342 2267
rect 6342 2215 6344 2267
rect 6288 2213 6344 2215
rect 6839 3551 6895 3607
rect 6703 2213 6759 2269
rect 6288 777 6344 779
rect 6288 725 6290 777
rect 6290 725 6342 777
rect 6342 725 6344 777
rect 6288 723 6344 725
rect 6567 723 6623 779
rect 12772 6434 12828 6436
rect 12772 6382 12774 6434
rect 12774 6382 12826 6434
rect 12826 6382 12828 6434
rect 12772 6380 12828 6382
<< metal3 >>
rect 38876 41201 38942 41204
rect 39379 41201 39445 41204
rect 38876 41199 39445 41201
rect 38876 41143 38881 41199
rect 38937 41143 39384 41199
rect 39440 41143 39445 41199
rect 38876 41141 39445 41143
rect 38876 41138 38942 41141
rect 39379 41138 39445 41141
rect 10994 40193 30885 40259
rect 10994 39871 30885 39937
rect 38604 39711 38670 39714
rect 39379 39711 39445 39714
rect 38604 39709 39445 39711
rect 38604 39653 38609 39709
rect 38665 39653 39384 39709
rect 39440 39653 39445 39709
rect 38604 39651 39445 39653
rect 38604 39648 38670 39651
rect 39379 39648 39445 39651
rect 10994 39033 30885 39099
rect 38740 38373 38806 38376
rect 39379 38373 39445 38376
rect 38740 38371 39445 38373
rect 10994 38259 30885 38325
rect 38740 38315 38745 38371
rect 38801 38315 39384 38371
rect 39440 38315 39445 38371
rect 38740 38313 39445 38315
rect 38740 38310 38806 38313
rect 39379 38310 39445 38313
rect 35058 38170 35124 38173
rect 20907 38168 35124 38170
rect 20907 38112 35063 38168
rect 35119 38112 35124 38168
rect 20907 38110 35124 38112
rect 35058 38107 35124 38110
rect 38876 37454 38942 37457
rect 32818 37452 38942 37454
rect 32818 37396 38881 37452
rect 38937 37396 38942 37452
rect 32818 37394 38942 37396
rect 38876 37391 38942 37394
rect 38604 37330 38670 37333
rect 32818 37328 38670 37330
rect 32818 37272 38609 37328
rect 38665 37272 38670 37328
rect 32818 37270 38670 37272
rect 38604 37267 38670 37270
rect 38740 37206 38806 37209
rect 32818 37204 38806 37206
rect 32818 37148 38745 37204
rect 38801 37148 38806 37204
rect 32818 37146 38806 37148
rect 38740 37143 38806 37146
rect 38604 37082 38670 37085
rect 32818 37080 38670 37082
rect 32818 37024 38609 37080
rect 38665 37024 38670 37080
rect 32818 37022 38670 37024
rect 38604 37019 38670 37022
rect 38604 36883 38670 36886
rect 39379 36883 39445 36886
rect 38604 36881 39445 36883
rect 38604 36825 38609 36881
rect 38665 36825 39384 36881
rect 39440 36825 39445 36881
rect 38604 36823 39445 36825
rect 38604 36820 38670 36823
rect 39379 36820 39445 36823
rect 10994 36262 32271 36328
rect 32895 35544 32961 35547
rect 32895 35542 45812 35544
rect 32895 35486 32900 35542
rect 32956 35486 45812 35542
rect 32895 35484 45812 35486
rect 32895 35481 32961 35484
rect 35182 35395 35248 35398
rect 22249 35393 35248 35395
rect 22249 35337 35187 35393
rect 35243 35337 35248 35393
rect 22249 35335 35248 35337
rect 35182 35332 35248 35335
rect 10994 34729 33505 34795
rect 38467 33768 38565 33866
rect 2290 14229 2388 14327
rect 2715 14229 2813 14327
rect 3094 14222 3192 14320
rect 3490 14222 3588 14320
rect 42140 14222 42238 14320
rect 42536 14222 42634 14320
rect 42915 14229 43013 14327
rect 43340 14229 43438 14327
rect 996 13432 1094 13530
rect 1392 13432 1490 13530
rect 2290 13439 2388 13537
rect 2715 13439 2813 13537
rect 3094 13432 3192 13530
rect 3490 13432 3588 13530
rect 42140 13432 42238 13530
rect 42536 13432 42634 13530
rect 42915 13439 43013 13537
rect 43340 13439 43438 13537
rect 44238 13432 44336 13530
rect 44634 13432 44732 13530
rect 2290 11859 2388 11957
rect 2715 11859 2813 11957
rect 3094 11852 3192 11950
rect 3490 11852 3588 11950
rect 42140 11852 42238 11950
rect 42536 11852 42634 11950
rect 42915 11859 43013 11957
rect 43340 11859 43438 11957
rect 996 11062 1094 11160
rect 1392 11062 1490 11160
rect 2290 11069 2388 11167
rect 2715 11069 2813 11167
rect 3094 11062 3192 11160
rect 3490 11062 3588 11160
rect 42140 11062 42238 11160
rect 42536 11062 42634 11160
rect 42915 11069 43013 11167
rect 43340 11069 43438 11167
rect 44238 11062 44336 11160
rect 44634 11062 44732 11160
rect 2290 9489 2388 9587
rect 2715 9489 2813 9587
rect 3094 9482 3192 9580
rect 3490 9482 3588 9580
rect 42140 9482 42238 9580
rect 42536 9482 42634 9580
rect 42915 9489 43013 9587
rect 43340 9489 43438 9587
rect 996 8692 1094 8790
rect 1392 8692 1490 8790
rect 2290 8699 2388 8797
rect 2715 8699 2813 8797
rect 3094 8692 3192 8790
rect 3490 8692 3588 8790
rect 42140 8692 42238 8790
rect 42536 8692 42634 8790
rect 42915 8699 43013 8797
rect 43340 8699 43438 8797
rect 44238 8692 44336 8790
rect 44634 8692 44732 8790
rect 7163 8106 7261 8204
rect 10994 7127 32881 7193
rect 10446 6587 10512 6590
rect 10446 6585 21937 6587
rect 10446 6529 10451 6585
rect 10507 6529 21937 6585
rect 10446 6527 21937 6529
rect 10446 6524 10512 6527
rect 12767 6438 12833 6441
rect 0 6436 12833 6438
rect 0 6380 12772 6436
rect 12828 6380 12833 6436
rect 0 6378 12833 6380
rect 12767 6375 12833 6378
rect 10994 5594 32271 5660
rect 6283 5099 6349 5102
rect 6562 5099 6628 5102
rect 6283 5097 6628 5099
rect 6283 5041 6288 5097
rect 6344 5041 6567 5097
rect 6623 5041 6628 5097
rect 6283 5039 6628 5041
rect 6283 5036 6349 5039
rect 6562 5036 6628 5039
rect 6562 4900 6628 4903
rect 6562 4898 10991 4900
rect 6562 4842 6567 4898
rect 6623 4842 10991 4898
rect 6562 4840 10991 4842
rect 6562 4837 6628 4840
rect 6834 4776 6900 4779
rect 6834 4774 10991 4776
rect 6834 4718 6839 4774
rect 6895 4718 10991 4774
rect 6834 4716 10991 4718
rect 6834 4713 6900 4716
rect 6698 4652 6764 4655
rect 6698 4650 10991 4652
rect 6698 4594 6703 4650
rect 6759 4594 10991 4650
rect 6698 4592 10991 4594
rect 6698 4589 6764 4592
rect 6562 4528 6628 4531
rect 6562 4526 10991 4528
rect 6562 4470 6567 4526
rect 6623 4470 10991 4526
rect 6562 4468 10991 4470
rect 6562 4465 6628 4468
rect 6283 3609 6349 3612
rect 6834 3609 6900 3612
rect 6283 3607 6900 3609
rect 6283 3551 6288 3607
rect 6344 3551 6839 3607
rect 6895 3551 6900 3607
rect 6283 3549 6900 3551
rect 6283 3546 6349 3549
rect 6834 3546 6900 3549
rect 10994 3378 30885 3444
rect 10994 2941 30885 3007
rect 10994 2609 30885 2675
rect 6283 2271 6349 2274
rect 6698 2271 6764 2274
rect 6283 2269 6764 2271
rect 6283 2213 6288 2269
rect 6344 2213 6703 2269
rect 6759 2213 6764 2269
rect 6283 2211 6764 2213
rect 6283 2208 6349 2211
rect 6698 2208 6764 2211
rect 10994 2117 30885 2183
rect 6283 781 6349 784
rect 6562 781 6628 784
rect 6283 779 6628 781
rect 6283 723 6288 779
rect 6344 723 6567 779
rect 6623 723 6628 779
rect 6283 721 6628 723
rect 6283 718 6349 721
rect 6562 718 6628 721
<< metal4 >>
rect 40011 36151 40077 41873
rect 41221 36102 41287 41922
rect 5022 8313 5088 33687
rect 5494 8313 5560 33687
rect 5926 8313 5992 33687
rect 6270 8313 6336 33687
rect 6694 8313 6760 33687
rect 7586 8283 7652 33689
rect 8011 8281 8077 33691
rect 8654 8313 8720 33659
rect 9902 8313 9968 33659
rect 11003 7506 11069 34416
rect 11413 7506 11479 34416
rect 34249 7506 34315 34416
rect 34659 7506 34725 34416
rect 35760 8313 35826 33659
rect 37008 8313 37074 33659
rect 37651 8281 37717 33691
rect 38076 8283 38142 33689
rect 38968 8313 39034 33687
rect 39392 8313 39458 33687
rect 39736 8313 39802 33687
rect 40168 8313 40234 33687
rect 40640 8313 40706 33687
rect 4441 0 4507 5820
rect 5651 49 5717 5771
use subbyte2_capped_replica_bitcell_array  subbyte2_capped_replica_bitcell_array_0
timestamp 1543373562
transform 1 0 10961 0 1 7506
box 0 0 23806 26910
use subbyte2_column_decoder  subbyte2_column_decoder_0
timestamp 1543373571
transform -1 0 41611 0 -1 41840
box 0 -82 2390 5738
use subbyte2_column_decoder  subbyte2_column_decoder_1
timestamp 1543373571
transform 1 0 4117 0 1 82
box 0 -82 2390 5738
use subbyte2_port_address  subbyte2_port_address_0
timestamp 1543373569
transform 1 0 0 0 1 8346
box 0 -490 10689 25345
use subbyte2_port_address_0  subbyte2_port_address_0_0
timestamp 1543373570
transform -1 0 45728 0 1 8346
box 0 -65 10689 25770
use subbyte2_port_data  subbyte2_port_data_0
timestamp 1543373570
transform 1 0 10961 0 -1 7506
box 0 252 21920 5669
use subbyte2_port_data_0  subbyte2_port_data_0_0
timestamp 1543373570
transform 1 0 10961 0 1 34416
box 0 252 22544 6218
<< labels >>
rlabel metal2 s 10465 82 10493 7506 4 p_en_bar0
port 3 nsew
rlabel metal2 s 10589 82 10617 7506 4 w_en0
port 5 nsew
rlabel metal2 s 7438 8033 7466 8061 4 wl_en0
port 7 nsew
rlabel metal2 s 35077 34416 35105 41924 4 s_en1
port 9 nsew
rlabel metal2 s 35201 34416 35229 41924 4 p_en_bar1
port 11 nsew
rlabel metal2 s 38262 33911 38290 33939 4 wl_en1
port 13 nsew
rlabel metal1 s 13103 1837 13163 1893 4 din0_0
port 15 nsew
rlabel metal1 s 15599 1837 15659 1893 4 din0_1
port 17 nsew
rlabel metal1 s 18095 1837 18155 1893 4 din0_2
port 19 nsew
rlabel metal1 s 20591 1837 20651 1893 4 din0_3
port 21 nsew
rlabel metal1 s 23087 1837 23147 1893 4 din0_4
port 23 nsew
rlabel metal1 s 25583 1837 25643 1893 4 din0_5
port 25 nsew
rlabel metal1 s 28079 1837 28139 1893 4 din0_6
port 27 nsew
rlabel metal1 s 30575 1837 30635 1893 4 din0_7
port 29 nsew
rlabel metal3 s 0 6378 12800 6438 4 rbl_bl_0_0
port 31 nsew
rlabel metal1 s 19 8346 47 14666 4 addr0_2
port 33 nsew
rlabel metal1 s 99 8346 127 14666 4 addr0_3
port 35 nsew
rlabel metal1 s 179 8346 207 14666 4 addr0_4
port 37 nsew
rlabel metal1 s 259 8346 287 14666 4 addr0_5
port 39 nsew
rlabel metal1 s 339 8346 367 14666 4 addr0_6
port 41 nsew
rlabel metal1 s 419 8346 447 14666 4 addr0_7
port 43 nsew
rlabel metal1 s 4232 722 4278 780 4 addr0_0
port 45 nsew
rlabel metal1 s 4356 2212 4402 2270 4 addr0_1
port 47 nsew
rlabel metal1 s 12984 40484 13030 40634 4 dout1_0
port 49 nsew
rlabel metal1 s 15480 40484 15526 40634 4 dout1_1
port 51 nsew
rlabel metal1 s 17976 40484 18022 40634 4 dout1_2
port 53 nsew
rlabel metal1 s 20472 40484 20518 40634 4 dout1_3
port 55 nsew
rlabel metal1 s 22968 40484 23014 40634 4 dout1_4
port 57 nsew
rlabel metal1 s 25464 40484 25510 40634 4 dout1_5
port 59 nsew
rlabel metal1 s 27960 40484 28006 40634 4 dout1_6
port 61 nsew
rlabel metal1 s 30456 40484 30502 40634 4 dout1_7
port 63 nsew
rlabel metal3 s 32928 35484 45812 35544 4 rbl_bl_1_1
port 65 nsew
rlabel metal1 s 45681 8346 45709 14666 4 addr1_2
port 67 nsew
rlabel metal1 s 45601 8346 45629 14666 4 addr1_3
port 69 nsew
rlabel metal1 s 45521 8346 45549 14666 4 addr1_4
port 71 nsew
rlabel metal1 s 45441 8346 45469 14666 4 addr1_5
port 73 nsew
rlabel metal1 s 45361 8346 45389 14666 4 addr1_6
port 75 nsew
rlabel metal1 s 45281 8346 45309 14666 4 addr1_7
port 77 nsew
rlabel metal1 s 41450 41142 41496 41200 4 addr1_0
port 79 nsew
rlabel metal1 s 41326 39652 41372 39710 4 addr1_1
port 81 nsew
rlabel metal3 s 3490 9482 3588 9580 4 vdd
port 83 nsew
rlabel metal3 s 42140 11062 42238 11160 4 vdd
port 83 nsew
rlabel metal4 s 5651 49 5717 5771 4 vdd
port 83 nsew
rlabel metal3 s 42915 11069 43013 11167 4 vdd
port 83 nsew
rlabel metal3 s 42915 11859 43013 11957 4 vdd
port 83 nsew
rlabel metal3 s 10994 2117 30885 2183 4 vdd
port 83 nsew
rlabel metal4 s 38968 8313 39034 33687 4 vdd
port 83 nsew
rlabel metal3 s 1392 13432 1490 13530 4 vdd
port 83 nsew
rlabel metal4 s 5494 8313 5560 33687 4 vdd
port 83 nsew
rlabel metal3 s 7163 8106 7261 8204 4 vdd
port 83 nsew
rlabel metal4 s 5926 8313 5992 33687 4 vdd
port 83 nsew
rlabel metal4 s 40168 8313 40234 33687 4 vdd
port 83 nsew
rlabel metal3 s 42915 8699 43013 8797 4 vdd
port 83 nsew
rlabel metal3 s 2715 9489 2813 9587 4 vdd
port 83 nsew
rlabel metal4 s 8011 8281 8077 33691 4 vdd
port 83 nsew
rlabel metal1 s 8019 7944 8069 8378 4 vdd
port 83 nsew
rlabel metal3 s 42915 13439 43013 13537 4 vdd
port 83 nsew
rlabel metal3 s 42140 8692 42238 8790 4 vdd
port 83 nsew
rlabel metal3 s 2715 11859 2813 11957 4 vdd
port 83 nsew
rlabel metal3 s 44238 11062 44336 11160 4 vdd
port 83 nsew
rlabel metal3 s 3490 11852 3588 11950 4 vdd
port 83 nsew
rlabel metal3 s 42915 14229 43013 14327 4 vdd
port 83 nsew
rlabel metal3 s 42140 14222 42238 14320 4 vdd
port 83 nsew
rlabel metal3 s 10994 39033 30885 39099 4 vdd
port 83 nsew
rlabel metal1 s 37659 33594 37709 34028 4 vdd
port 83 nsew
rlabel metal3 s 2715 13439 2813 13537 4 vdd
port 83 nsew
rlabel metal4 s 34659 7506 34725 34416 4 vdd
port 83 nsew
rlabel metal3 s 42140 11852 42238 11950 4 vdd
port 83 nsew
rlabel metal4 s 39736 8313 39802 33687 4 vdd
port 83 nsew
rlabel metal1 s 35779 33626 35807 34021 4 vdd
port 83 nsew
rlabel metal3 s 2715 11069 2813 11167 4 vdd
port 83 nsew
rlabel metal3 s 10994 34729 33505 34795 4 vdd
port 83 nsew
rlabel metal3 s 1392 8692 1490 8790 4 vdd
port 83 nsew
rlabel metal3 s 1392 11062 1490 11160 4 vdd
port 83 nsew
rlabel metal3 s 10994 39871 30885 39937 4 vdd
port 83 nsew
rlabel metal4 s 9902 8313 9968 33659 4 vdd
port 83 nsew
rlabel metal3 s 44238 13432 44336 13530 4 vdd
port 83 nsew
rlabel metal4 s 6694 8313 6760 33687 4 vdd
port 83 nsew
rlabel metal3 s 3490 8692 3588 8790 4 vdd
port 83 nsew
rlabel metal3 s 42915 9489 43013 9587 4 vdd
port 83 nsew
rlabel metal3 s 3490 11062 3588 11160 4 vdd
port 83 nsew
rlabel metal1 s 9921 7951 9949 8346 4 vdd
port 83 nsew
rlabel metal4 s 40011 36151 40077 41873 4 vdd
port 83 nsew
rlabel metal3 s 3490 13432 3588 13530 4 vdd
port 83 nsew
rlabel metal3 s 2715 8699 2813 8797 4 vdd
port 83 nsew
rlabel metal3 s 38467 33768 38565 33866 4 vdd
port 83 nsew
rlabel metal4 s 35760 8313 35826 33659 4 vdd
port 83 nsew
rlabel metal3 s 42140 13432 42238 13530 4 vdd
port 83 nsew
rlabel metal3 s 2715 14229 2813 14327 4 vdd
port 83 nsew
rlabel metal3 s 44238 8692 44336 8790 4 vdd
port 83 nsew
rlabel metal3 s 10994 2941 30885 3007 4 vdd
port 83 nsew
rlabel metal3 s 42140 9482 42238 9580 4 vdd
port 83 nsew
rlabel metal4 s 37651 8281 37717 33691 4 vdd
port 83 nsew
rlabel metal3 s 10994 7127 32881 7193 4 vdd
port 83 nsew
rlabel metal3 s 3490 14222 3588 14320 4 vdd
port 83 nsew
rlabel metal4 s 11003 7506 11069 34416 4 vdd
port 83 nsew
rlabel metal3 s 3094 14222 3192 14320 4 gnd
port 85 nsew
rlabel metal3 s 10994 40193 30885 40259 4 gnd
port 85 nsew
rlabel metal3 s 3094 9482 3192 9580 4 gnd
port 85 nsew
rlabel metal3 s 42536 8692 42634 8790 4 gnd
port 85 nsew
rlabel metal3 s 2290 14229 2388 14327 4 gnd
port 85 nsew
rlabel metal3 s 42536 13432 42634 13530 4 gnd
port 85 nsew
rlabel metal4 s 4441 0 4507 5820 4 gnd
port 85 nsew
rlabel metal3 s 2290 13439 2388 13537 4 gnd
port 85 nsew
rlabel metal3 s 3094 11062 3192 11160 4 gnd
port 85 nsew
rlabel metal3 s 42536 9482 42634 9580 4 gnd
port 85 nsew
rlabel metal3 s 43340 11069 43438 11167 4 gnd
port 85 nsew
rlabel metal3 s 44634 8692 44732 8790 4 gnd
port 85 nsew
rlabel metal4 s 5022 8313 5088 33687 4 gnd
port 85 nsew
rlabel metal3 s 2290 11069 2388 11167 4 gnd
port 85 nsew
rlabel metal4 s 39392 8313 39458 33687 4 gnd
port 85 nsew
rlabel metal4 s 6270 8313 6336 33687 4 gnd
port 85 nsew
rlabel metal3 s 10994 36262 32271 36328 4 gnd
port 85 nsew
rlabel metal4 s 37008 8313 37074 33659 4 gnd
port 85 nsew
rlabel metal4 s 40640 8313 40706 33687 4 gnd
port 85 nsew
rlabel metal4 s 8654 8313 8720 33659 4 gnd
port 85 nsew
rlabel metal4 s 34249 7506 34315 34416 4 gnd
port 85 nsew
rlabel metal3 s 10994 3378 30885 3444 4 gnd
port 85 nsew
rlabel metal3 s 42536 14222 42634 14320 4 gnd
port 85 nsew
rlabel metal4 s 11413 7506 11479 34416 4 gnd
port 85 nsew
rlabel metal3 s 10994 38259 30885 38325 4 gnd
port 85 nsew
rlabel metal3 s 42536 11062 42634 11160 4 gnd
port 85 nsew
rlabel metal3 s 2290 9489 2388 9587 4 gnd
port 85 nsew
rlabel metal3 s 3094 8692 3192 8790 4 gnd
port 85 nsew
rlabel metal4 s 7586 8283 7652 33689 4 gnd
port 85 nsew
rlabel metal3 s 42536 11852 42634 11950 4 gnd
port 85 nsew
rlabel metal3 s 44634 11062 44732 11160 4 gnd
port 85 nsew
rlabel metal3 s 44634 13432 44732 13530 4 gnd
port 85 nsew
rlabel metal3 s 10994 5594 32271 5660 4 gnd
port 85 nsew
rlabel metal4 s 41221 36102 41287 41922 4 gnd
port 85 nsew
rlabel metal3 s 2290 8699 2388 8797 4 gnd
port 85 nsew
rlabel metal3 s 996 13432 1094 13530 4 gnd
port 85 nsew
rlabel metal3 s 996 8692 1094 8790 4 gnd
port 85 nsew
rlabel metal3 s 43340 14229 43438 14327 4 gnd
port 85 nsew
rlabel metal3 s 10994 2609 30885 2675 4 gnd
port 85 nsew
rlabel metal3 s 43340 11859 43438 11957 4 gnd
port 85 nsew
rlabel metal3 s 996 11062 1094 11160 4 gnd
port 85 nsew
rlabel metal3 s 3094 11852 3192 11950 4 gnd
port 85 nsew
rlabel metal3 s 3094 13432 3192 13530 4 gnd
port 85 nsew
rlabel metal3 s 2290 11859 2388 11957 4 gnd
port 85 nsew
rlabel metal3 s 43340 13439 43438 13537 4 gnd
port 85 nsew
rlabel metal3 s 43340 8699 43438 8797 4 gnd
port 85 nsew
rlabel metal3 s 43340 9489 43438 9587 4 gnd
port 85 nsew
rlabel metal4 s 38076 8283 38142 33689 4 gnd
port 85 nsew
<< properties >>
string FIXED_BBOX 0 0 45812 41842
<< end >>
