* NGSPICE file created from subbyte2.ext - technology: sky130A

.subckt subbyte2_pnand2_0 A B Z vdd gnd
X0 a_144_51# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.259p pd=2.18u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd B Z vdd sky130_fd_pr__pfet_01v8 ad=0.672p pd=5.68u as=0.392p ps=2.94u w=1.12u l=0.15u
X2 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z B a_144_51# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt subbyte2_pinv_3 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=2.4696p pd=16.38u as=2.4696p ps=16.38u w=1.68u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=2.94p pd=18.94u as=2.94p ps=18.94u w=2u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X8 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X9 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X10 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X11 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pdriver_0 A Z vdd gnd
Xsubbyte2_pinv_3_0 A Z vdd gnd subbyte2_pinv_3
.ends

.subckt subbyte2_pnand2 A B Z vdd w_n36_679# gnd
X0 a_144_51# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.259p pd=2.18u as=0.222p ps=2.08u w=0.74u l=0.15u
X1 vdd B Z w_n36_679# sky130_fd_pr__pfet_01v8 ad=0.672p pd=5.68u as=0.392p ps=2.94u w=1.12u l=0.15u
X2 Z A vdd w_n36_679# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z B a_144_51# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt subbyte2_pand2_0 A B Z gnd vdd
Xsubbyte2_pdriver_0_0 subbyte2_pnand2_0/Z Z vdd gnd subbyte2_pdriver_0
Xsubbyte2_pnand2_0 A B subbyte2_pnand2_0/Z vdd vdd gnd subbyte2_pnand2
.ends

.subckt subbyte2_pinv_10 A Z vdd gnd
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=4.68p pd=28.68u as=5.1p ps=33.1u w=2u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=4.68p pd=28.68u as=5.1p ps=33.1u w=2u l=0.15u
X2 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pinv_9 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.9828p pd=6.6u as=1.2474p ps=9.54u w=1.26u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=1.56p pd=9.56u as=1.98p ps=13.98u w=2u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt subbyte2_pdriver_2 A Z vdd gnd
Xsubbyte2_pinv_10_0 subbyte2_pinv_9_0/Z Z vdd gnd subbyte2_pinv_10
Xsubbyte2_pinv_9_0 A subbyte2_pinv_9_0/Z vdd gnd subbyte2_pinv_9
.ends

.subckt subbyte2_pinv_13 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt subbyte2_delay_chain in out vdd gnd
Xsubbyte2_pinv_13_8 subbyte2_pinv_13_9/Z subbyte2_pinv_13_8/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_13 subbyte2_pinv_13_9/A subbyte2_pinv_13_13/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_24 subbyte2_pinv_13_29/Z subbyte2_pinv_13_24/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_35 subbyte2_pinv_13_39/Z subbyte2_pinv_13_35/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_9 subbyte2_pinv_13_9/A subbyte2_pinv_13_9/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_14 subbyte2_pinv_13_19/Z subbyte2_pinv_13_9/A vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_25 subbyte2_pinv_13_29/Z subbyte2_pinv_13_25/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_36 subbyte2_pinv_13_39/Z subbyte2_pinv_13_36/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_15 subbyte2_pinv_13_19/Z subbyte2_pinv_13_15/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_26 subbyte2_pinv_13_29/Z subbyte2_pinv_13_26/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_37 subbyte2_pinv_13_39/Z subbyte2_pinv_13_37/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_16 subbyte2_pinv_13_19/Z subbyte2_pinv_13_16/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_27 subbyte2_pinv_13_29/Z subbyte2_pinv_13_27/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_38 subbyte2_pinv_13_39/Z subbyte2_pinv_13_38/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_17 subbyte2_pinv_13_19/Z subbyte2_pinv_13_17/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_28 subbyte2_pinv_13_29/Z subbyte2_pinv_13_28/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_39 subbyte2_pinv_13_44/Z subbyte2_pinv_13_39/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_18 subbyte2_pinv_13_19/Z subbyte2_pinv_13_18/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_29 subbyte2_pinv_13_34/Z subbyte2_pinv_13_29/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_19 subbyte2_pinv_13_24/Z subbyte2_pinv_13_19/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_0 out subbyte2_pinv_13_0/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_1 out subbyte2_pinv_13_1/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_2 out subbyte2_pinv_13_2/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_40 subbyte2_pinv_13_44/Z subbyte2_pinv_13_40/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_3 out subbyte2_pinv_13_3/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_30 subbyte2_pinv_13_34/Z subbyte2_pinv_13_30/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_41 subbyte2_pinv_13_44/Z subbyte2_pinv_13_41/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_4 subbyte2_pinv_13_9/Z out vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_20 subbyte2_pinv_13_24/Z subbyte2_pinv_13_20/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_31 subbyte2_pinv_13_34/Z subbyte2_pinv_13_31/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_42 subbyte2_pinv_13_44/Z subbyte2_pinv_13_42/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_5 subbyte2_pinv_13_9/Z subbyte2_pinv_13_5/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_6 subbyte2_pinv_13_9/Z subbyte2_pinv_13_6/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_10 subbyte2_pinv_13_9/A subbyte2_pinv_13_10/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_11 subbyte2_pinv_13_9/A subbyte2_pinv_13_11/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_21 subbyte2_pinv_13_24/Z subbyte2_pinv_13_21/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_22 subbyte2_pinv_13_24/Z subbyte2_pinv_13_22/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_32 subbyte2_pinv_13_34/Z subbyte2_pinv_13_32/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_33 subbyte2_pinv_13_34/Z subbyte2_pinv_13_33/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_43 subbyte2_pinv_13_44/Z subbyte2_pinv_13_43/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_44 in subbyte2_pinv_13_44/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_7 subbyte2_pinv_13_9/Z subbyte2_pinv_13_7/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_12 subbyte2_pinv_13_9/A subbyte2_pinv_13_12/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_23 subbyte2_pinv_13_24/Z subbyte2_pinv_13_23/Z vdd gnd subbyte2_pinv_13
Xsubbyte2_pinv_13_34 subbyte2_pinv_13_39/Z subbyte2_pinv_13_34/Z vdd gnd subbyte2_pinv_13
.ends

.subckt subbyte2_pinv_0 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt subbyte2_pinv_6 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=1.1592p pd=8.1u as=1.1592p ps=8.1u w=1.68u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=1.1592p pd=8.1u as=1.1592p ps=8.1u w=1.68u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
.ends

.subckt subbyte2_pinv_7 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=2.34p pd=14.34u as=2.76p ps=18.76u w=2u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=2.34p pd=14.34u as=2.76p ps=18.76u w=2u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pinv A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt subbyte2_pdriver_5 A Z gnd vdd
Xsubbyte2_pinv_6_0 subbyte2_pinv_0/Z subbyte2_pinv_7_0/A vdd gnd subbyte2_pinv_6
Xsubbyte2_pinv_7_0 subbyte2_pinv_7_0/A Z vdd gnd subbyte2_pinv_7
Xsubbyte2_pinv_0 subbyte2_pinv_1/Z subbyte2_pinv_0/Z vdd gnd subbyte2_pinv
Xsubbyte2_pinv_1 A subbyte2_pinv_1/Z vdd gnd subbyte2_pinv
.ends

.subckt subbyte2_pinv_8 A Z vdd gnd
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=7.02p pd=43.02u as=7.44p ps=47.44u w=2u l=0.15u
X1 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X2 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=7.02p pd=43.02u as=7.44p ps=47.44u w=2u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X18 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X19 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X20 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X21 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X22 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X23 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X24 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X25 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X26 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X27 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X28 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X29 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X30 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X31 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X32 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X33 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X34 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X35 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pdriver_1 A Z gnd vdd
Xsubbyte2_pinv_8_0 subbyte2_pinv_8_0/A Z vdd gnd subbyte2_pinv_8
Xsubbyte2_pinv_6_0 subbyte2_pinv_0/Z subbyte2_pinv_7_0/A vdd gnd subbyte2_pinv_6
Xsubbyte2_pinv_7_0 subbyte2_pinv_7_0/A subbyte2_pinv_8_0/A vdd gnd subbyte2_pinv_7
Xsubbyte2_pinv_0 subbyte2_pinv_1/Z subbyte2_pinv_0/Z vdd gnd subbyte2_pinv
Xsubbyte2_pinv_2 A subbyte2_pinv_2/Z vdd gnd subbyte2_pinv
Xsubbyte2_pinv_1 subbyte2_pinv_2/Z subbyte2_pinv_1/Z vdd gnd subbyte2_pinv
.ends

.subckt subbyte2_pinv_12 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=1.8144p pd=12.24u as=1.8144p ps=12.24u w=1.68u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=2.16p pd=14.16u as=2.16p ps=14.16u w=2u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X8 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X9 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pdriver_4 A Z vdd gnd
Xsubbyte2_pinv_12_0 A Z vdd gnd subbyte2_pinv_12
.ends

.subckt subbyte2_pnand3 A B C Z vdd w_n36_679# gnd
X0 Z C vdd w_n36_679# sky130_fd_pr__pfet_01v8 ad=0.728p pd=5.78u as=0.728p ps=5.78u w=1.12u l=0.15u
X1 a_144_51# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.259p pd=2.18u as=0.222p ps=2.08u w=0.74u l=0.15u
X2 vdd B Z w_n36_679# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X3 Z A vdd w_n36_679# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X4 Z C a_244_51# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0.259p ps=2.18u w=0.74u l=0.15u
X5 a_244_51# B a_144_51# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt subbyte2_pand3_0 A B C Z vdd gnd
Xsubbyte2_pdriver_4_0 subbyte2_pnand3_0/Z Z vdd gnd subbyte2_pdriver_4
Xsubbyte2_pnand3_0 A B C subbyte2_pnand3_0/Z vdd vdd gnd subbyte2_pnand3
.ends

.subckt subbyte2_pinv_2 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=1.1592p pd=8.1u as=1.1592p ps=8.1u w=1.68u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X2 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=1.1592p pd=8.1u as=1.1592p ps=8.1u w=1.68u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68u l=0.15u
.ends

.subckt sky130_fd_bd_sram__openram_dff D Q gnd clk vdd QN
X0 vdd a_28_102# a_389_712# vdd sky130_fd_pr__pfet_01v8 ad=3.315p pd=26.21u as=0.63p ps=6.42u w=3u l=0.15u
X1 a_47_611# clk a_197_712# vdd sky130_fd_pr__pfet_01v8 ad=1.35p pd=6.9u as=0.63p ps=6.42u w=3u l=0.15u
X2 a_239_76# clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0.795p pd=6.53u as=0p ps=0u w=3u l=0.15u
X3 a_197_712# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X4 QN clk a_547_102# gnd sky130_fd_pr__nfet_01v8 ad=0.45p pd=2.9u as=0.21p ps=2.42u w=1u l=0.15u
X5 gnd Q a_739_102# gnd sky130_fd_pr__nfet_01v8 ad=1.105p pd=10.21u as=0.21p ps=2.42u w=1u l=0.15u
X6 Q QN gnd gnd sky130_fd_pr__nfet_01v8 ad=0.265p pd=2.53u as=0p ps=0u w=1u l=0.15u
X7 a_389_712# a_239_76# a_47_611# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X8 vdd a_47_611# a_28_102# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0.795p ps=6.53u w=3u l=0.15u
X9 a_547_712# a_28_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63p pd=6.42u as=0p ps=0u w=3u l=0.15u
X10 a_739_712# clk QN vdd sky130_fd_pr__pfet_01v8 ad=0.63p pd=6.42u as=1.35p ps=6.9u w=3u l=0.15u
X11 gnd a_28_102# a_389_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.21p ps=2.42u w=1u l=0.15u
X12 a_47_611# a_239_76# a_197_102# gnd sky130_fd_pr__nfet_01v8 ad=0.45p pd=2.9u as=0.21p ps=2.42u w=1u l=0.15u
X13 a_239_76# clk gnd gnd sky130_fd_pr__nfet_01v8 ad=0.265p pd=2.53u as=0p ps=0u w=1u l=0.15u
X14 a_197_102# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1u l=0.15u
X15 a_389_102# clk a_47_611# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1u l=0.15u
X16 gnd a_47_611# a_28_102# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.265p ps=2.53u w=1u l=0.15u
X17 a_547_102# a_28_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1u l=0.15u
X18 a_739_102# a_239_76# QN gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1u l=0.15u
X19 vdd Q a_739_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X20 QN a_239_76# a_547_712# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X21 Q QN vdd vdd sky130_fd_pr__pfet_01v8 ad=0.795p pd=6.53u as=0p ps=0u w=3u l=0.15u
.ends

.subckt subbyte2_pinv_1 A Z vdd gnd
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.2886p pd=2.26u as=0.444p ps=4.16u w=0.74u l=0.15u
X1 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.74u l=0.15u
X2 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0.756p pd=6.24u as=0.4914p ps=3.3u w=1.26u l=0.15u
X3 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
.ends

.subckt subbyte2_dff_buf_0 Q Qb clk vdd gnd D
Xsubbyte2_pinv_2_0 Qb Q vdd gnd subbyte2_pinv_2
Xsky130_fd_bd_sram__openram_dff_0 D subbyte2_pinv_1_0/A gnd clk vdd sky130_fd_bd_sram__openram_dff_0/QN
+ sky130_fd_bd_sram__openram_dff
Xsubbyte2_pinv_1_0 subbyte2_pinv_1_0/A Qb vdd gnd subbyte2_pinv_1
.ends

.subckt subbyte2_dff_buf_array dout_0 clk dout_bar_0 vdd din_0 gnd
Xsubbyte2_dff_buf_0_0 dout_0 dout_bar_0 clk vdd gnd din_0 subbyte2_dff_buf_0
.ends

.subckt subbyte2_control_logic_r clk rbl_bl s_en p_en_bar wl_en clk_buf vdd_uq1 csb
+ vdd gnd vdd_uq0
Xsubbyte2_pnand2_0_0 subbyte2_pand2_0_0/Z subbyte2_pand3_0_0/A subbyte2_pnand2_0_0/Z
+ vdd_uq1 gnd subbyte2_pnand2_0
Xsubbyte2_pand2_0_1 subbyte2_pinv_0_0/Z subbyte2_pand3_0_0/C subbyte2_pand3_0_0/B
+ gnd vdd_uq1 subbyte2_pand2_0
Xsubbyte2_pdriver_2_0 subbyte2_pand3_0_0/B wl_en vdd_uq1 gnd subbyte2_pdriver_2
Xsubbyte2_delay_chain_0 rbl_bl subbyte2_pand3_0_0/A vdd_uq0 gnd subbyte2_delay_chain
Xsubbyte2_pinv_0_0 clk_buf subbyte2_pinv_0_0/Z vdd_uq1 gnd subbyte2_pinv_0
Xsubbyte2_pdriver_5_0 subbyte2_pnand2_0_0/Z p_en_bar gnd vdd_uq1 subbyte2_pdriver_5
Xsubbyte2_pdriver_1_0 clk clk_buf gnd vdd_uq1 subbyte2_pdriver_1
Xsubbyte2_pand3_0_0 subbyte2_pand3_0_0/A subbyte2_pand3_0_0/B subbyte2_pand3_0_0/C
+ s_en vdd_uq1 gnd subbyte2_pand3_0
Xsubbyte2_dff_buf_array_0 subbyte2_dff_buf_array_0/dout_0 clk_buf subbyte2_pand3_0_0/C
+ vdd csb gnd subbyte2_dff_buf_array
Xsubbyte2_pand2_0_0 clk_buf subbyte2_pand3_0_0/C subbyte2_pand2_0_0/Z gnd vdd_uq1
+ subbyte2_pand2_0
.ends

.subckt subbyte2_pinv_11 A Z vdd gnd
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=3.72p pd=23.72u as=3.72p ps=23.72u w=2u l=0.15u
X1 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=3.72p pd=23.72u as=3.72p ps=23.72u w=2u l=0.15u
X2 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X3 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X4 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X5 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X6 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X7 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X8 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X9 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X10 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X11 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X12 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X13 Z A gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X14 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X15 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X16 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
X17 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u
.ends

.subckt subbyte2_pdriver_3 A Z vdd gnd
Xsubbyte2_pinv_11_0 A Z vdd gnd subbyte2_pinv_11
.ends

.subckt subbyte2_pand3 A B C Z vdd gnd
Xsubbyte2_pdriver_3_0 subbyte2_pnand3_0/Z Z vdd gnd subbyte2_pdriver_3
Xsubbyte2_pnand3_0 A B C subbyte2_pnand3_0/Z vdd vdd gnd subbyte2_pnand3
.ends

.subckt subbyte2_control_logic_w clk rbl_bl w_en p_en_bar wl_en clk_buf vdd_uq1 csb
+ gnd vdd vdd_uq0
Xsubbyte2_pnand2_0_0 subbyte2_pand2_0_0/Z subbyte2_pinv_0_0/A subbyte2_pnand2_0_0/Z
+ vdd_uq1 gnd subbyte2_pnand2_0
Xsubbyte2_pand2_0_1 subbyte2_pinv_0_1/Z subbyte2_pand3_0/A subbyte2_pand3_0/C gnd
+ vdd_uq1 subbyte2_pand2_0
Xsubbyte2_pdriver_2_0 subbyte2_pand3_0/C wl_en vdd_uq1 gnd subbyte2_pdriver_2
Xsubbyte2_delay_chain_0 rbl_bl subbyte2_pinv_0_0/A vdd_uq0 gnd subbyte2_delay_chain
Xsubbyte2_pinv_0_0 subbyte2_pinv_0_0/A subbyte2_pand3_0/B vdd_uq1 gnd subbyte2_pinv_0
Xsubbyte2_pinv_0_1 clk_buf subbyte2_pinv_0_1/Z vdd_uq1 gnd subbyte2_pinv_0
Xsubbyte2_pdriver_5_0 subbyte2_pnand2_0_0/Z p_en_bar gnd vdd_uq1 subbyte2_pdriver_5
Xsubbyte2_pdriver_1_0 clk clk_buf gnd vdd_uq1 subbyte2_pdriver_1
Xsubbyte2_dff_buf_array_0 subbyte2_dff_buf_array_0/dout_0 clk_buf subbyte2_pand3_0/A
+ vdd csb gnd subbyte2_dff_buf_array
Xsubbyte2_pand3_0 subbyte2_pand3_0/A subbyte2_pand3_0/B subbyte2_pand3_0/C w_en vdd_uq1
+ gnd subbyte2_pand3
Xsubbyte2_pand2_0_0 clk_buf subbyte2_pand3_0/A subbyte2_pand2_0_0/Z gnd vdd_uq1 subbyte2_pand2_0
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell gnd bl0 br0 bl1 br1 wl0 wl1 vdd a_38_n79#
+ a_400_n79#
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=1.0032p pd=13.14u as=0.0504p ps=0.9u w=0.21u l=0.08u
X1 a_38_133# wl0 a_38_133# vdd sky130_fd_pr__special_pfet_pass ad=0.035p pd=0.78u as=0p ps=0u w=0.07u l=0.15u
X2 a_16_183# wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0.3088p pd=4.43u as=0.0504p ps=0.9u w=0.21u l=0.15u
X3 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X4 a_16_183# a_38_133# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.2768p ps=4u w=0.21u l=0.15u
X5 a_16_183# wl1 a_16_183# vdd sky130_fd_pr__special_pfet_pass ad=0.035p pd=0.78u as=0p ps=0u w=0.07u l=0.15u
X6 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0.3463p pd=4.93u as=0p ps=0u w=0.21u l=0.15u
X7 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X8 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.08u
X9 a_38_133# a_16_183# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X10 br0 wl0 a_16_183# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.105p ps=1.84u w=0.21u l=0.15u
X11 gnd a_38_133# a_16_183# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X12 a_38_133# a_16_183# vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0.0364p ps=0.8u w=0.14u l=0.15u
X13 vdd a_38_133# a_16_183# vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=0.14u l=0.15u
X14 bl0 wl0 a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.105p ps=1.84u w=0.21u l=0.15u
X15 gnd a_16_183# a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
.ends

.subckt subbyte2_bitcell_array bl_1_12 br_0_19 bl_1_23 wl_0_2 wl_0_15 wl_0_16 wl_0_17
+ wl_0_26 wl_0_37 wl_0_38 wl_0_48 wl_0_49 wl_1_53 wl_1_62 wl_1_63 vdd_uq222 vdd_uq318
+ vdd_uq446 vdd_uq478 vdd_uq510 vdd_uq638 vdd_uq670 vdd_uq830 vdd_uq990 sky130_fd_bd_sram__openram_dp_cell_447/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1407/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_0/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_960/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1024/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_576/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_895/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1536/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1855/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_767/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1471/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2047/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1279/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_320/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1984/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1023/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1535/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_320/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_768/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1472/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_192/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1152/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_319/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1471/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_127/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1279/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1536/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_64/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_448/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_767/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1408/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_831/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1983/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1727/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_511/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_128/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_896/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1856/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_575/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1599/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_640/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_832/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1984/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1600/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_0/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_383/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1024/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1343/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_639/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1343/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_576/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1280/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1600/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1472/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_639/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1791/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1087/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1407/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1344/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_768/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1728/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1791/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_512/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_831/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1088/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_63/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1408/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_255/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_383/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1215/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_703/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1855/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_960/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_640/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1792/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1920/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_384/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1344/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1663/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_447/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1151/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1599/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_64/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1919/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1087/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_384/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_704/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1856/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1792/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_959/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1919/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1215/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_448/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1152/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_703/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_2047/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_127/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_895/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_832/a_38_n79#
+ wl_0_25 sky130_fd_bd_sram__openram_dp_cell_1216/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_256/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_575/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1216/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_191/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1535/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_511/a_400_n79# wl_1_8 sky130_fd_bd_sram__openram_dp_cell_959/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1663/a_400_n79# wl_0_53 sky130_fd_bd_sram__openram_dp_cell_896/a_400_n79#
+ wl_0_8 sky130_fd_bd_sram__openram_dp_cell_1920/a_400_n79# wl_1_16 wl_0_63 wl_1_7
+ sky130_fd_bd_sram__openram_dp_cell_1664/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1983/a_38_n79#
+ wl_0_7 wl_0_62 sky130_fd_bd_sram__openram_dp_cell_255/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1088/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_1727/a_400_n79# wl_1_44 wl_1_35 sky130_fd_bd_sram__openram_dp_cell_192/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_512/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1664/a_400_n79#
+ wl_0_44 wl_0_29 bl_0_21 sky130_fd_bd_sram__openram_dp_cell_191/a_38_n79# bl_0_1
+ wl_0_35 br_1_31 wl_1_28 br_0_18 bl_0_4 wl_1_11 vdd_uq94 vdd_uq734 wl_0_58 bl_1_20
+ wl_1_2 wl_1_57 br_0_25 br_0_5 bl_0_11 br_0_1 bl_0_7 br_1_17 wl_1_22 sky130_fd_bd_sram__openram_dp_cell_1151/a_38_n79#
+ wl_1_13 bl_1_26 br_1_20 bl_1_6 br_0_24 vdd_uq542 bl_0_10 wl_0_5 br_0_4 wl_0_60 wl_1_54
+ br_1_23 bl_1_29 br_1_3 bl_1_9 bl_0_17 vdd_uq958 bl_0_31 br_0_7 bl_0_30 wl_1_42 wl_0_46
+ wl_1_19 wl_1_33 vdd_uq190 sky130_fd_bd_sram__openram_dp_cell_319/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_1023/a_400_n79#
+ wl_1_45 br_0_31 wl_1_24 br_1_30 br_1_10 vdd_uq862 wl_0_20 vdd_uq350 wl_0_28 bl_0_24
+ br_0_14 wl_1_36 wl_0_11 bl_1_16 br_1_26 wl_0_19 br_1_6 bl_0_0 bl_0_20 wl_1_27 bl_1_19
+ wl_1_18 wl_1_10 br_1_29 br_1_9 bl_1_15 wl_0_57 wl_1_9 wl_1_1 wl_0_40 vdd_uq894 br_1_16
+ wl_1_0 wl_1_48 br_1_13 wl_1_56 wl_0_31 bl_0_2 br_0_17 bl_0_23 bl_0_3 br_1_12 wl_1_55
+ wl_1_39 vdd_uq766 vdd_uq99 wl_0_22 br_0_21 bl_0_27 wl_1_46 wl_1_30 wl_1_38 wl_1_25
+ wl_0_13 bl_0_26 br_0_20 bl_0_6 br_1_11 wl_1_37 wl_1_21 bl_0_25 wl_1_29 bl_1_2 bl_1_22
+ bl_1_18 wl_1_4 wl_1_12 wl_0_51 sky130_fd_bd_sram__openram_dp_cell_704/a_38_n79#
+ bl_1_0 wl_1_59 wl_1_3 bl_0_5 bl_1_1 bl_1_21 vdd_uq574 vdd_uq702 wl_0_30 br_0_27
+ bl_0_13 wl_1_50 sky130_fd_bd_sram__openram_dp_cell_256/a_400_n79# br_1_15 wl_0_21
+ wl_0_54 br_0_23 br_0_3 wl_1_41 bl_0_29 bl_0_9 br_1_19 bl_1_25 bl_1_5 vdd wl_1_47
+ br_0_0 br_1_22 bl_1_28 br_1_2 bl_1_8 wl_0_4 br_1_14 bl_1_24 wl_0_12 bl_0_28 wl_1_20
+ br_1_18 bl_1_4 wl_1_15 wl_0_3 br_0_22 wl_0_42 wl_0_50 bl_1_3 bl_0_8 wl_1_58 wl_0_33
+ vdd_uq606 wl_0_41 br_0_2 wl_0_45 vdd_uq62 wl_1_49 wl_0_24 wl_0_32 br_0_30 br_0_10
+ wl_0_36 wl_1_32 br_0_28 vdd_uq254 wl_1_40 bl_1_27 sky130_fd_bd_sram__openram_dp_cell_1728/a_400_n79#
+ wl_0_23 bl_0_16 br_0_6 bl_0_12 br_0_26 wl_0_27 wl_1_23 bl_0_14 vdd_uq382 wl_1_31
+ br_1_5 br_1_25 wl_0_6 br_1_21 wl_1_26 wl_0_14 bl_0_19 wl_1_6 wl_0_18 br_0_8 wl_1_14
+ bl_1_11 wl_0_10 wl_0_61 wl_1_17 br_1_1 bl_1_7 br_0_29 br_0_9 bl_0_15 wl_1_61 wl_0_9
+ wl_1_5 wl_0_1 wl_0_52 br_1_0 sky130_fd_bd_sram__openram_dp_cell_128/a_38_n79# br_0_16
+ wl_1_52 wl_0_0 wl_1_60 sky130_fd_bd_sram__openram_dp_cell_1280/a_38_n79# vdd_uq414
+ wl_0_56 wl_0_43 br_0_13 br_1_27 vdd_uq999 wl_0_59 sky130_fd_bd_sram__openram_dp_cell_63/a_38_n79#
+ br_0_12 wl_1_43 vdd_uq286 wl_0_55 br_1_28 bl_1_17 wl_0_39 wl_1_51 bl_1_14 br_1_8
+ vdd_uq926 br_1_24 br_1_4 wl_0_47 bl_1_10 wl_0_34 bl_1_30 bl_0_22 bl_0_18 br_1_7
+ bl_1_13 gnd br_0_15 vdd_uq798 br_0_11 wl_1_34 bl_1_31 vdd_uq158
Xsky130_fd_bd_sram__openram_dp_cell_262 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_57
+ wl_1_57 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_251 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_4
+ wl_1_4 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_240 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_15
+ wl_1_15 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_295 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_24
+ wl_1_24 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_284 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_35
+ wl_1_35 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_273 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_46
+ wl_1_46 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1409 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_62 wl_1_62
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_806 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_25
+ wl_1_25 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1921 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_62 wl_1_62
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_839 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_56
+ wl_1_56 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1910 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_9 wl_1_9
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_828 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_3
+ wl_1_3 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_817 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_14
+ wl_1_14 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1987 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_60 wl_1_60
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1932 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_51 wl_1_51
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1998 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_49 wl_1_49
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1976 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_7 wl_1_7
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1965 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_18 wl_1_18
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1954 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_29 wl_1_29
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1943 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_40 wl_1_40
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1217 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_62
+ wl_1_62 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1206 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_9
+ wl_1_9 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1228 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_51
+ wl_1_51 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1239 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_40
+ wl_1_40 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_647 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_56
+ wl_1_56 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_636 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_3
+ wl_1_3 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_625 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_14
+ wl_1_14 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_614 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_25
+ wl_1_25 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_603 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_36
+ wl_1_36 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1740 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_51 wl_1_51
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1762 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_29 wl_1_29
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_669 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_34
+ wl_1_34 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1751 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_40 wl_1_40
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_658 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_45
+ wl_1_45 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1795 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_60 wl_1_60
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1784 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_7 wl_1_7
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1773 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_18 wl_1_18
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1025 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_62
+ wl_1_62 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1036 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_51
+ wl_1_51 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1014 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_9
+ wl_1_9 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1003 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_20
+ wl_1_20 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1058 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_29
+ wl_1_29 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1047 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_40
+ wl_1_40 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1069 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_18
+ wl_1_18 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_455 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_56
+ wl_1_56 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_400 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_47
+ wl_1_47 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_444 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_3
+ wl_1_3 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_499 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_12
+ wl_1_12 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_433 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_14
+ wl_1_14 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_488 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_23
+ wl_1_23 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_422 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_25
+ wl_1_25 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_477 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_34
+ wl_1_34 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_411 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_36
+ wl_1_36 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_466 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_45
+ wl_1_45 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1592 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_7 wl_1_7
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1581 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_18 wl_1_18
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1570 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_29 wl_1_29
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_263 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_56
+ wl_1_56 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_252 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_3
+ wl_1_3 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_241 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_14
+ wl_1_14 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_296 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_23
+ wl_1_23 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_230 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_25
+ wl_1_25 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_285 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_34
+ wl_1_34 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_274 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_45
+ wl_1_45 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_829 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_2
+ wl_1_2 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_818 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_13
+ wl_1_13 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_807 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_24
+ wl_1_24 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1922 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_61 wl_1_61
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1933 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_50 wl_1_50
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1911 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_8 wl_1_8
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1900 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_19 wl_1_19
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1955 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_28 wl_1_28
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1944 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_39 wl_1_39
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1988 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_59 wl_1_59
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1977 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_6 wl_1_6
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1966 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_17 wl_1_17
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1999 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_48 wl_1_48
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1218 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_61
+ wl_1_61 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1229 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_50
+ wl_1_50 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1207 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_8
+ wl_1_8 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_648 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_55
+ wl_1_55 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_637 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_2
+ wl_1_2 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_626 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_13
+ wl_1_13 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_615 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_24
+ wl_1_24 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_604 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_35
+ wl_1_35 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_659 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_44
+ wl_1_44 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1730 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_61 wl_1_61
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1796 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_59 wl_1_59
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1741 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_50 wl_1_50
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1785 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_6 wl_1_6
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1774 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_17 wl_1_17
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1763 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_28 wl_1_28
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1752 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_39 wl_1_39
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1026 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_61
+ wl_1_61 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1037 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_50
+ wl_1_50 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1015 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_8
+ wl_1_8 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1004 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_19
+ wl_1_19 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1059 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_28
+ wl_1_28 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1048 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_39
+ wl_1_39 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_456 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_55
+ wl_1_55 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_445 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_2
+ wl_1_2 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_434 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_13
+ wl_1_13 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_489 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_22
+ wl_1_22 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_423 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_24
+ wl_1_24 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_478 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_33
+ wl_1_33 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_412 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_35
+ wl_1_35 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_467 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_44
+ wl_1_44 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_401 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_46
+ wl_1_46 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1593 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_6 wl_1_6
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1582 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_17 wl_1_17
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1571 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_28 wl_1_28
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1560 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_39 wl_1_39
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_990 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_33
+ wl_1_33 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_231 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_24
+ wl_1_24 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_220 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_35
+ wl_1_35 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_264 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_55
+ wl_1_55 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_253 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_2
+ wl_1_2 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_242 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_13
+ wl_1_13 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_297 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_22
+ wl_1_22 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_286 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_33
+ wl_1_33 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_275 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_44
+ wl_1_44 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1390 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_17
+ wl_1_17 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_819 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_12
+ wl_1_12 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_808 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_23
+ wl_1_23 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1923 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_60 wl_1_60
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1934 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_49 wl_1_49
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1912 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_7 wl_1_7
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1978 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_5 wl_1_5
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1967 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_16 wl_1_16
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1901 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_18 wl_1_18
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1956 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_27 wl_1_27
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1945 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_38 wl_1_38
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1989 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_58 wl_1_58
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1219 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_60
+ wl_1_60 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1208 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_7
+ wl_1_7 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_649 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_54
+ wl_1_54 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_638 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_1
+ wl_1_1 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_627 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_12
+ wl_1_12 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_616 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_23
+ wl_1_23 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_605 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_34
+ wl_1_34 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1731 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_60 wl_1_60
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1797 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_58 wl_1_58
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1742 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_49 wl_1_49
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1720 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_7 wl_1_7
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1786 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_5 wl_1_5
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1775 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_16 wl_1_16
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1764 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_27 wl_1_27
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1753 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_38 wl_1_38
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1027 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_60
+ wl_1_60 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1038 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_49
+ wl_1_49 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1016 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_7
+ wl_1_7 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1005 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_18
+ wl_1_18 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1049 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_38
+ wl_1_38 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_413 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_34
+ wl_1_34 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_402 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_45
+ wl_1_45 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_457 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_54
+ wl_1_54 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_446 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_1
+ wl_1_1 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_435 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_12
+ wl_1_12 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_424 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_23
+ wl_1_23 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_479 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_32
+ wl_1_32 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_468 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_43
+ wl_1_43 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1550 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_49 wl_1_49
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1594 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_5 wl_1_5
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1583 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_16 wl_1_16
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1572 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_27 wl_1_27
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1561 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_38 wl_1_38
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_991 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_32
+ wl_1_32 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_980 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_43
+ wl_1_43 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_265 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_54
+ wl_1_54 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_254 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_1
+ wl_1_1 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_243 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_12
+ wl_1_12 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_232 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_23
+ wl_1_23 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_221 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_34
+ wl_1_34 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_210 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_45
+ wl_1_45 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_298 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_21
+ wl_1_21 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1380 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_27
+ wl_1_27 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_287 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_32
+ wl_1_32 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_276 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_43
+ wl_1_43 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1391 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_16
+ wl_1_16 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_809 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_22
+ wl_1_22 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1924 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_59 wl_1_59
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1913 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_6 wl_1_6
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1979 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_4 wl_1_4
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1968 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_15 wl_1_15
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1902 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_17 wl_1_17
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1957 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_26 wl_1_26
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1946 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_37 wl_1_37
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1935 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_48 wl_1_48
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1209 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_6
+ wl_1_6 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1721 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_6 wl_1_6
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_639 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_0
+ wl_1_0 vdd_uq318 sky130_fd_bd_sram__openram_dp_cell_639/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_639/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_628 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_11
+ wl_1_11 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1710 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_17 wl_1_17
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_617 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_22
+ wl_1_22 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_606 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_33
+ wl_1_33 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1732 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_59 wl_1_59
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1798 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_57 wl_1_57
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1787 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_4 wl_1_4
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1776 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_15 wl_1_15
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1765 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_26 wl_1_26
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1754 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_37 wl_1_37
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1743 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_48 wl_1_48
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1006 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_17
+ wl_1_17 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1028 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_59
+ wl_1_59 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1017 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_6
+ wl_1_6 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1039 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_48
+ wl_1_48 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_447 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_0
+ wl_1_0 vdd_uq222 sky130_fd_bd_sram__openram_dp_cell_447/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_447/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_436 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_11
+ wl_1_11 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_425 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_22
+ wl_1_22 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_414 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_33
+ wl_1_33 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_403 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_44
+ wl_1_44 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1540 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_59 wl_1_59
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_458 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_53
+ wl_1_53 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1562 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_37 wl_1_37
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_469 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_42
+ wl_1_42 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1551 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_48 wl_1_48
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1595 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_4 wl_1_4
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1584 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_15 wl_1_15
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1573 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_26 wl_1_26
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_970 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_53
+ wl_1_53 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_992 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_31
+ wl_1_31 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_981 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_42
+ wl_1_42 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_200 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_55
+ wl_1_55 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_266 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_53
+ wl_1_53 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_255 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_0
+ wl_1_0 vdd_uq99 sky130_fd_bd_sram__openram_dp_cell_255/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_255/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_244 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_11
+ wl_1_11 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_233 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_22
+ wl_1_22 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_288 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_31
+ wl_1_31 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_222 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_33
+ wl_1_33 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_277 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_42
+ wl_1_42 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_211 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_44
+ wl_1_44 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1392 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_15
+ wl_1_15 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_299 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_20
+ wl_1_20 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1381 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_26
+ wl_1_26 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1370 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_37
+ wl_1_37 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_90 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_37
+ wl_1_37 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1903 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_16 wl_1_16
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1925 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_58 wl_1_58
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1914 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_5 wl_1_5
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1969 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_14 wl_1_14
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1958 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_25 wl_1_25
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1947 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_36 wl_1_36
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1936 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_47 wl_1_47
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_629 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_10
+ wl_1_10 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_618 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_21
+ wl_1_21 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_607 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_32
+ wl_1_32 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1733 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_58 wl_1_58
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1722 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_5 wl_1_5
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1711 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_16 wl_1_16
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1700 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_27 wl_1_27
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1744 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_47 wl_1_47
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1799 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_56 wl_1_56
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1788 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_3 wl_1_3
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1777 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_14 wl_1_14
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1766 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_25 wl_1_25
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1755 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_36 wl_1_36
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1029 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_58
+ wl_1_58 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1018 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_5
+ wl_1_5 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1007 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_16
+ wl_1_16 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_448 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_63
+ wl_1_63 vdd_uq254 sky130_fd_bd_sram__openram_dp_cell_448/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_448/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_459 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_52
+ wl_1_52 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_437 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_10
+ wl_1_10 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_426 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_21
+ wl_1_21 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_415 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_32
+ wl_1_32 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_404 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_43
+ wl_1_43 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1541 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_58 wl_1_58
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1530 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_5 wl_1_5
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1596 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_3 wl_1_3
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1585 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_14 wl_1_14
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1574 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_25 wl_1_25
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1563 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_36 wl_1_36
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1552 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_47 wl_1_47
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_960 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_63
+ wl_1_63 vdd_uq510 sky130_fd_bd_sram__openram_dp_cell_960/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_960/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_971 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_52
+ wl_1_52 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_993 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_30
+ wl_1_30 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_982 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_41
+ wl_1_41 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_256 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_63
+ wl_1_63 vdd_uq158 sky130_fd_bd_sram__openram_dp_cell_256/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_256/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_201 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_54
+ wl_1_54 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_267 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_52
+ wl_1_52 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_245 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_10
+ wl_1_10 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_234 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_21
+ wl_1_21 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_289 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_30
+ wl_1_30 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_223 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_32
+ wl_1_32 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_278 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_41
+ wl_1_41 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_212 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_43
+ wl_1_43 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1393 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_14
+ wl_1_14 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1382 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_25
+ wl_1_25 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1371 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_36
+ wl_1_36 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1360 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_47
+ wl_1_47 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_790 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_41
+ wl_1_41 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_80 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_47
+ wl_1_47 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_91 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_36
+ wl_1_36 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1190 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_25
+ wl_1_25 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1926 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_57 wl_1_57
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1915 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_4 wl_1_4
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1904 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_15 wl_1_15
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1937 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_46 wl_1_46
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1959 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_24 wl_1_24
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1948 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_35 wl_1_35
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_619 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_20
+ wl_1_20 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_608 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_31
+ wl_1_31 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1734 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_57 wl_1_57
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1723 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_4 wl_1_4
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1778 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_13 wl_1_13
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1712 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_15 wl_1_15
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1767 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_24 wl_1_24
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1701 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_26 wl_1_26
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1756 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_35 wl_1_35
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1745 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_46 wl_1_46
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1789 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_2 wl_1_2
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1019 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_4
+ wl_1_4 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1008 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_15
+ wl_1_15 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_449 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_62
+ wl_1_62 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_438 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_9
+ wl_1_9 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_427 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_20
+ wl_1_20 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_416 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_31
+ wl_1_31 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_405 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_42
+ wl_1_42 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1542 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_57 wl_1_57
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1531 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_4 wl_1_4
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1597 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_2 wl_1_2
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1586 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_13 wl_1_13
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1520 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_15 wl_1_15
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1575 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_24 wl_1_24
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1564 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_35 wl_1_35
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1553 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_46 wl_1_46
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_961 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_62
+ wl_1_62 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_972 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_51
+ wl_1_51 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_950 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_9
+ wl_1_9 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_994 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_29
+ wl_1_29 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_983 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_40
+ wl_1_40 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_202 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_53
+ wl_1_53 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_213 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_42
+ wl_1_42 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_257 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_62
+ wl_1_62 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_268 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_51
+ wl_1_51 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_246 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_9
+ wl_1_9 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2040 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_7 wl_1_7
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_235 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_20
+ wl_1_20 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_224 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_31
+ wl_1_31 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_279 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_40
+ wl_1_40 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1350 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_57
+ wl_1_57 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1394 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_13
+ wl_1_13 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1383 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_24
+ wl_1_24 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1372 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_35
+ wl_1_35 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1361 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_46
+ wl_1_46 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_780 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_51
+ wl_1_51 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_791 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_40
+ wl_1_40 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_70 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_57
+ wl_1_57 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_92 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_35
+ wl_1_35 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_81 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_46
+ wl_1_46 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1191 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_24
+ wl_1_24 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1180 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_35
+ wl_1_35 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1927 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_56 wl_1_56
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1916 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_3 wl_1_3
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1905 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_14 wl_1_14
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1949 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_34 wl_1_34
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1938 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_45 wl_1_45
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_609 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_30
+ wl_1_30 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1735 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_56 wl_1_56
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1779 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_12 wl_1_12
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1724 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_3 wl_1_3
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1713 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_14 wl_1_14
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1768 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_23 wl_1_23
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1702 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_25 wl_1_25
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1757 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_34 wl_1_34
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1746 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_45 wl_1_45
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1009 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_14
+ wl_1_14 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_439 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_8
+ wl_1_8 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_428 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_19
+ wl_1_19 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1510 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_25 wl_1_25
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_417 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_30
+ wl_1_30 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_406 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_41
+ wl_1_41 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1543 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_56 wl_1_56
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1587 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_12 wl_1_12
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1532 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_3 wl_1_3
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1598 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_1 wl_1_1
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1521 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_14 wl_1_14
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1576 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_23 wl_1_23
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1565 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_34 wl_1_34
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1554 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_45 wl_1_45
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_951 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_8
+ wl_1_8 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_940 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_19
+ wl_1_19 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_962 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_61
+ wl_1_61 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_973 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_50
+ wl_1_50 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_995 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_28
+ wl_1_28 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_984 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_39
+ wl_1_39 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_203 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_52
+ wl_1_52 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_247 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_8
+ wl_1_8 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_236 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_19
+ wl_1_19 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_225 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_30
+ wl_1_30 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_214 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_41
+ wl_1_41 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_258 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_61
+ wl_1_61 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1351 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_56
+ wl_1_56 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_269 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_50
+ wl_1_50 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2041 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_6 wl_1_6
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1340 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_3
+ wl_1_3 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2030 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_17 wl_1_17
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1362 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_45
+ wl_1_45 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1395 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_12
+ wl_1_12 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1384 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_23
+ wl_1_23 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1373 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_34
+ wl_1_34 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_770 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_61
+ wl_1_61 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_781 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_50
+ wl_1_50 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_792 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_39
+ wl_1_39 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_71 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_56
+ wl_1_56 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_60 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_3
+ wl_1_3 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1192 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_23
+ wl_1_23 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1181 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_34
+ wl_1_34 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_93 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_34
+ wl_1_34 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1170 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_45
+ wl_1_45 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_82 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_45
+ wl_1_45 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1928 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_55 wl_1_55
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1917 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_2 wl_1_2
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1906 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_13 wl_1_13
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1939 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_44 wl_1_44
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1703 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_24 wl_1_24
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1736 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_55 wl_1_55
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1725 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_2 wl_1_2
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1714 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_13 wl_1_13
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1769 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_22 wl_1_22
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1758 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_33 wl_1_33
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1747 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_44 wl_1_44
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_429 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_18
+ wl_1_18 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_418 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_29
+ wl_1_29 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_407 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_40
+ wl_1_40 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1544 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_55 wl_1_55
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1533 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_2 wl_1_2
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1522 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_13 wl_1_13
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1511 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_24 wl_1_24
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1500 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_35 wl_1_35
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1588 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_11 wl_1_11
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1599 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_0 wl_1_0
+ vdd_uq798 sky130_fd_bd_sram__openram_dp_cell_1599/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1599/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1577 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_22 wl_1_22
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1566 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_33 wl_1_33
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1555 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_44 wl_1_44
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_963 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_60
+ wl_1_60 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_974 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_49
+ wl_1_49 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_952 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_7
+ wl_1_7 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_941 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_18
+ wl_1_18 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_930 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_29
+ wl_1_29 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_985 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_38
+ wl_1_38 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_996 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_27
+ wl_1_27 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_259 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_60
+ wl_1_60 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_204 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_51
+ wl_1_51 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_248 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_7
+ wl_1_7 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_237 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_18
+ wl_1_18 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_226 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_29
+ wl_1_29 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_215 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_40
+ wl_1_40 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1352 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_55
+ wl_1_55 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1396 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_11
+ wl_1_11 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2042 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_5 wl_1_5
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1341 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_2
+ wl_1_2 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1330 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_13
+ wl_1_13 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2031 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_16 wl_1_16
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1385 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_22
+ wl_1_22 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2020 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_27 wl_1_27
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1374 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_33
+ wl_1_33 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1363 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_44
+ wl_1_44 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_0 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_63
+ wl_1_63 vdd sky130_fd_bd_sram__openram_dp_cell_0/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_0/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_771 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_60
+ wl_1_60 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_782 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_49
+ wl_1_49 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_760 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_7
+ wl_1_7 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_793 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_38
+ wl_1_38 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_50 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_13
+ wl_1_13 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_72 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_55
+ wl_1_55 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1160 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_55
+ wl_1_55 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_61 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_2
+ wl_1_2 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1193 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_22
+ wl_1_22 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1182 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_33
+ wl_1_33 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_94 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_33
+ wl_1_33 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1171 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_44
+ wl_1_44 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_83 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_44
+ wl_1_44 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_590 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_49
+ wl_1_49 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1929 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_54 wl_1_54
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1907 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_12 wl_1_12
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1918 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_1 wl_1_1
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1715 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_12 wl_1_12
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1726 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_1 wl_1_1
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1704 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_23 wl_1_23
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1737 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_54 wl_1_54
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1759 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_32 wl_1_32
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1748 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_43 wl_1_43
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_419 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_28
+ wl_1_28 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_408 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_39
+ wl_1_39 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1545 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_54 wl_1_54
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1523 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_12 wl_1_12
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1534 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_1 wl_1_1
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1578 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_21 wl_1_21
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1512 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_23 wl_1_23
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1567 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_32 wl_1_32
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1501 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_34 wl_1_34
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1556 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_43 wl_1_43
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1589 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_10 wl_1_10
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_964 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_59
+ wl_1_59 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_975 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_48
+ wl_1_48 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_953 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_6
+ wl_1_6 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_942 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_17
+ wl_1_17 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_997 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_26
+ wl_1_26 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_931 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_28
+ wl_1_28 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_986 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_37
+ wl_1_37 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_920 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_39
+ wl_1_39 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_205 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_50
+ wl_1_50 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_249 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_6
+ wl_1_6 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_238 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_17
+ wl_1_17 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2021 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_26 wl_1_26
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_227 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_28
+ wl_1_28 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2010 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_37 wl_1_37
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_216 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_39
+ wl_1_39 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1353 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_54
+ wl_1_54 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1331 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_12
+ wl_1_12 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1397 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_10
+ wl_1_10 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2043 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_4 wl_1_4
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1342 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_1
+ wl_1_1 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2032 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_15 wl_1_15
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1386 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_21
+ wl_1_21 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1320 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_23
+ wl_1_23 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1375 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_32
+ wl_1_32 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1364 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_43
+ wl_1_43 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_62
+ wl_1_62 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_772 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_59
+ wl_1_59 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_783 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_48
+ wl_1_48 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_761 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_6
+ wl_1_6 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_750 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_17
+ wl_1_17 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_794 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_37
+ wl_1_37 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_73 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_54
+ wl_1_54 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_62 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_1
+ wl_1_1 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_51 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_12
+ wl_1_12 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_40 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_23
+ wl_1_23 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_84 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_43
+ wl_1_43 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1161 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_54
+ wl_1_54 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1150 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_1
+ wl_1_1 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1194 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_21
+ wl_1_21 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1183 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_32
+ wl_1_32 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_95 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_32
+ wl_1_32 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1172 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_43
+ wl_1_43 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_580 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_59
+ wl_1_59 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_591 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_48
+ wl_1_48 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1908 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_11 wl_1_11
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1919 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_0 wl_1_0
+ vdd_uq958 sky130_fd_bd_sram__openram_dp_cell_1919/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1919/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1738 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_53 wl_1_53
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1716 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_11 wl_1_11
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1727 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_0 wl_1_0
+ vdd_uq862 sky130_fd_bd_sram__openram_dp_cell_1727/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1727/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1705 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_22 wl_1_22
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1749 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_42 wl_1_42
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_409 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_38
+ wl_1_38 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1546 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_53 wl_1_53
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1524 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_11 wl_1_11
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1535 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_0 wl_1_0
+ vdd_uq766 sky130_fd_bd_sram__openram_dp_cell_1535/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1535/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1579 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_20 wl_1_20
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1513 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_22 wl_1_22
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1568 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_31 wl_1_31
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1502 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_33 wl_1_33
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1557 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_42 wl_1_42
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_965 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_58
+ wl_1_58 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_910 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_49
+ wl_1_49 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_976 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_47
+ wl_1_47 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_954 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_5
+ wl_1_5 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_943 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_16
+ wl_1_16 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_998 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_25
+ wl_1_25 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_932 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_27
+ wl_1_27 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_987 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_36
+ wl_1_36 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_921 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_38
+ wl_1_38 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_206 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_49
+ wl_1_49 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2044 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_3 wl_1_3
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2033 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_14 wl_1_14
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_239 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_16
+ wl_1_16 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2022 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_25 wl_1_25
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_228 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_27
+ wl_1_27 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1310 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_33
+ wl_1_33 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2011 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_36 wl_1_36
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_217 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_38
+ wl_1_38 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2000 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_47 wl_1_47
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1354 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_53
+ wl_1_53 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1332 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_11
+ wl_1_11 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1398 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_9
+ wl_1_9 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1343 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_0
+ wl_1_0 vdd_uq670 sky130_fd_bd_sram__openram_dp_cell_1343/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1343/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1387 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_20
+ wl_1_20 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1321 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_22
+ wl_1_22 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1376 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_31
+ wl_1_31 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1365 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_42
+ wl_1_42 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_61
+ wl_1_61 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_751 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_16
+ wl_1_16 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_740 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_27
+ wl_1_27 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_773 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_58
+ wl_1_58 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_784 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_47
+ wl_1_47 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_762 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_5
+ wl_1_5 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_795 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_36
+ wl_1_36 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_74 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_53
+ wl_1_53 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1140 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_11
+ wl_1_11 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1151 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_0
+ wl_1_0 vdd_uq574 sky130_fd_bd_sram__openram_dp_cell_1151/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1151/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_63 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_0
+ wl_1_0 vdd sky130_fd_bd_sram__openram_dp_cell_63/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_63/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_52 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_11
+ wl_1_11 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_41 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_22
+ wl_1_22 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_96 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_31
+ wl_1_31 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_30 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_33
+ wl_1_33 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_85 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_42
+ wl_1_42 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1162 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_53
+ wl_1_53 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1195 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_20
+ wl_1_20 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1184 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_31
+ wl_1_31 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1173 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_42
+ wl_1_42 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_581 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_58
+ wl_1_58 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_592 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_47
+ wl_1_47 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_570 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_5
+ wl_1_5 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1909 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_10 wl_1_10
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1728 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_63 wl_1_63
+ vdd_uq894 sky130_fd_bd_sram__openram_dp_cell_1728/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1728/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1739 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_52 wl_1_52
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1717 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_10 wl_1_10
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1706 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_21 wl_1_21
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1536 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_63 wl_1_63
+ vdd_uq798 sky130_fd_bd_sram__openram_dp_cell_1536/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1536/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1547 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_52 wl_1_52
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1525 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_10 wl_1_10
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1514 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_21 wl_1_21
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1569 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_30 wl_1_30
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1503 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_32 wl_1_32
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1558 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_41 wl_1_41
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_900 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_59
+ wl_1_59 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_911 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_48
+ wl_1_48 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_933 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_26
+ wl_1_26 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_922 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_37
+ wl_1_37 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_966 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_57
+ wl_1_57 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_955 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_4
+ wl_1_4 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_944 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_15
+ wl_1_15 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_999 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_24
+ wl_1_24 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_988 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_35
+ wl_1_35 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_977 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_46
+ wl_1_46 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_207 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_48
+ wl_1_48 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_229 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_26
+ wl_1_26 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_218 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_37
+ wl_1_37 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1344 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_63
+ wl_1_63 vdd_uq702 sky130_fd_bd_sram__openram_dp_cell_1344/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1344/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1333 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_10
+ wl_1_10 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2045 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_2 wl_1_2
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2034 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_13 wl_1_13
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1322 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_21
+ wl_1_21 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2023 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_24 wl_1_24
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1311 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_32
+ wl_1_32 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2012 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_35 wl_1_35
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1300 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_43
+ wl_1_43 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2001 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_46 wl_1_46
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1355 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_52
+ wl_1_52 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1399 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_8
+ wl_1_8 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1388 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_19
+ wl_1_19 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1377 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_30
+ wl_1_30 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1366 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_41
+ wl_1_41 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_3 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_60
+ wl_1_60 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_774 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_57
+ wl_1_57 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_763 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_4
+ wl_1_4 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_752 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_15
+ wl_1_15 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_741 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_26
+ wl_1_26 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_730 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_37
+ wl_1_37 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_796 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_35
+ wl_1_35 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_785 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_46
+ wl_1_46 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_64 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_63
+ wl_1_63 vdd_uq62 sky130_fd_bd_sram__openram_dp_cell_64/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_64/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1152 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_63
+ wl_1_63 vdd_uq606 sky130_fd_bd_sram__openram_dp_cell_1152/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1152/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_75 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_52
+ wl_1_52 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1163 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_52
+ wl_1_52 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_53 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_10
+ wl_1_10 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1141 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_10
+ wl_1_10 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1130 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_21
+ wl_1_21 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_42 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_21
+ wl_1_21 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1185 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_30
+ wl_1_30 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_97 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_30
+ wl_1_30 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_31 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_32
+ wl_1_32 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1174 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_41
+ wl_1_41 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_86 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_41
+ wl_1_41 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_20 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_43
+ wl_1_43 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1196 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_19
+ wl_1_19 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_582 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_57
+ wl_1_57 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_571 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_4
+ wl_1_4 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_560 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_15
+ wl_1_15 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_593 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_46
+ wl_1_46 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_390 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_57
+ wl_1_57 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1729 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_62 wl_1_62
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1718 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_9 wl_1_9
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1707 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_20 wl_1_20
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1526 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_9 wl_1_9
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1515 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_20 wl_1_20
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1504 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_31 wl_1_31
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1537 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_62 wl_1_62
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1548 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_51 wl_1_51
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1559 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_40 wl_1_40
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_901 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_58
+ wl_1_58 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_967 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_56
+ wl_1_56 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_912 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_47
+ wl_1_47 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_956 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_3
+ wl_1_3 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_945 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_14
+ wl_1_14 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_934 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_25
+ wl_1_25 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_923 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_36
+ wl_1_36 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_989 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_34
+ wl_1_34 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_978 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_45
+ wl_1_45 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_208 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_47
+ wl_1_47 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_219 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_36
+ wl_1_36 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1345 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_62
+ wl_1_62 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1356 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_51
+ wl_1_51 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2035 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_12 wl_1_12
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1334 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_9
+ wl_1_9 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2046 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_1 wl_1_1
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1323 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_20
+ wl_1_20 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2024 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_23 wl_1_23
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1312 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_31
+ wl_1_31 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2013 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_34 wl_1_34
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1367 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_40
+ wl_1_40 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1301 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_42
+ wl_1_42 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2002 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_45 wl_1_45
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1389 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_18
+ wl_1_18 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1378 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_29
+ wl_1_29 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_4 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_59
+ wl_1_59 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_775 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_56
+ wl_1_56 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_720 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_47
+ wl_1_47 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_764 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_3
+ wl_1_3 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_753 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_14
+ wl_1_14 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_742 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_25
+ wl_1_25 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_797 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_34
+ wl_1_34 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_731 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_36
+ wl_1_36 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_786 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_45
+ wl_1_45 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1890 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_29 wl_1_29
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_10 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_53
+ wl_1_53 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_32 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_31
+ wl_1_31 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_21 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_42
+ wl_1_42 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_65 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_62
+ wl_1_62 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1153 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_62
+ wl_1_62 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_76 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_51
+ wl_1_51 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1164 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_51
+ wl_1_51 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_54 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_9
+ wl_1_9 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1142 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_9
+ wl_1_9 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1197 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_18
+ wl_1_18 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1131 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_20
+ wl_1_20 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_43 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_20
+ wl_1_20 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1186 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_29
+ wl_1_29 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_98 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_29
+ wl_1_29 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1120 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_31
+ wl_1_31 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1175 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_40
+ wl_1_40 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_87 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_40
+ wl_1_40 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_583 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_56
+ wl_1_56 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_572 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_3
+ wl_1_3 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_561 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_14
+ wl_1_14 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_550 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_25
+ wl_1_25 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_594 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_45
+ wl_1_45 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_391 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_56
+ wl_1_56 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_380 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_3
+ wl_1_3 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1708 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_19 wl_1_19
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1719 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_8 wl_1_8
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1538 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_61 wl_1_61
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1549 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_50 wl_1_50
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1527 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_8 wl_1_8
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1516 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_19 wl_1_19
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1505 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_30 wl_1_30
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_902 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_57
+ wl_1_57 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_968 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_55
+ wl_1_55 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_957 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_2
+ wl_1_2 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_946 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_13
+ wl_1_13 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_935 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_24
+ wl_1_24 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_924 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_35
+ wl_1_35 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_979 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_44
+ wl_1_44 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_913 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_46
+ wl_1_46 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2003 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_44 wl_1_44
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_209 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_46
+ wl_1_46 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1346 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_61
+ wl_1_61 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1357 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_50
+ wl_1_50 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2036 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_11 wl_1_11
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1335 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_8
+ wl_1_8 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2047 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_0 wl_1_0
+ vdd_uq999 sky130_fd_bd_sram__openram_dp_cell_2047/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_2047/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1324 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_19
+ wl_1_19 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2025 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_22 wl_1_22
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1379 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_28
+ wl_1_28 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1313 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_30
+ wl_1_30 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2014 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_33 wl_1_33
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1368 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_39
+ wl_1_39 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1302 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_41
+ wl_1_41 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_5 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_58
+ wl_1_58 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_710 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_57
+ wl_1_57 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_776 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_55
+ wl_1_55 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_765 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_2
+ wl_1_2 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_754 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_13
+ wl_1_13 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_743 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_24
+ wl_1_24 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_798 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_33
+ wl_1_33 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_732 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_35
+ wl_1_35 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_787 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_44
+ wl_1_44 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_721 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_46
+ wl_1_46 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1891 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_28 wl_1_28
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1880 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_39 wl_1_39
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_66 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_61
+ wl_1_61 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_11 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_52
+ wl_1_52 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_55 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_8
+ wl_1_8 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_44 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_19
+ wl_1_19 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_33 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_30
+ wl_1_30 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1110 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_41
+ wl_1_41 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_22 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_41
+ wl_1_41 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1154 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_61
+ wl_1_61 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_77 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_50
+ wl_1_50 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1165 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_50
+ wl_1_50 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1143 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_8
+ wl_1_8 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1198 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_17
+ wl_1_17 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1132 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_19
+ wl_1_19 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1187 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_28
+ wl_1_28 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_99 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_28
+ wl_1_28 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1121 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_30
+ wl_1_30 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1176 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_39
+ wl_1_39 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_88 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_39
+ wl_1_39 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_540 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_35
+ wl_1_35 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_584 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_55
+ wl_1_55 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_573 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_2
+ wl_1_2 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_562 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_13
+ wl_1_13 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_551 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_24
+ wl_1_24 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_595 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_44
+ wl_1_44 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_392 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_55
+ wl_1_55 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_381 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_2
+ wl_1_2 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_370 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_13
+ wl_1_13 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1709 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_18 wl_1_18
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1539 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_60 wl_1_60
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1528 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_7 wl_1_7
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1517 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_18 wl_1_18
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1506 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_29 wl_1_29
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_903 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_56
+ wl_1_56 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_969 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_54
+ wl_1_54 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_958 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_1
+ wl_1_1 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_947 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_12
+ wl_1_12 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_936 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_23
+ wl_1_23 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_925 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_34
+ wl_1_34 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_914 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_45
+ wl_1_45 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2037 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_10 wl_1_10
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2026 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_21 wl_1_21
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2015 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_32 wl_1_32
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2004 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_43 wl_1_43
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1347 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_60
+ wl_1_60 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1358 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_49
+ wl_1_49 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1336 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_7
+ wl_1_7 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1325 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_18
+ wl_1_18 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1314 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_29
+ wl_1_29 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1369 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_38
+ wl_1_38 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1303 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_40
+ wl_1_40 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_6 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_57
+ wl_1_57 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_711 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_56
+ wl_1_56 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_700 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_3
+ wl_1_3 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_733 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_34
+ wl_1_34 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_722 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_45
+ wl_1_45 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_777 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_54
+ wl_1_54 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_766 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_1
+ wl_1_1 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_755 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_12
+ wl_1_12 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_744 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_23
+ wl_1_23 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_799 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_32
+ wl_1_32 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_788 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_43
+ wl_1_43 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1870 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_49 wl_1_49
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1892 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_27 wl_1_27
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1881 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_38 wl_1_38
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_67 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_60
+ wl_1_60 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_12 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_51
+ wl_1_51 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1100 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_51
+ wl_1_51 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_78 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_49
+ wl_1_49 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_56 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_7
+ wl_1_7 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1133 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_18
+ wl_1_18 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_45 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_18
+ wl_1_18 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1122 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_29
+ wl_1_29 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_34 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_29
+ wl_1_29 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_89 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_38
+ wl_1_38 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1111 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_40
+ wl_1_40 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_23 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_40
+ wl_1_40 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1155 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_60
+ wl_1_60 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1166 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_49
+ wl_1_49 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1144 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_7
+ wl_1_7 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1199 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_16
+ wl_1_16 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1188 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_27
+ wl_1_27 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1177 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_38
+ wl_1_38 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_574 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_1
+ wl_1_1 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_563 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_12
+ wl_1_12 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_552 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_23
+ wl_1_23 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_541 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_34
+ wl_1_34 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_530 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_45
+ wl_1_45 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_585 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_54
+ wl_1_54 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_596 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_43
+ wl_1_43 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_393 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_54
+ wl_1_54 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_382 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_1
+ wl_1_1 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_371 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_12
+ wl_1_12 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_360 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_23
+ wl_1_23 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_190 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_1
+ wl_1_1 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1529 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_6 wl_1_6
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1518 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_17 wl_1_17
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1507 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_28 wl_1_28
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_904 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_55
+ wl_1_55 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_915 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_44
+ wl_1_44 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_959 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_0
+ wl_1_0 vdd_uq478 sky130_fd_bd_sram__openram_dp_cell_959/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_959/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_948 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_11
+ wl_1_11 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_937 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_22
+ wl_1_22 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_926 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_33
+ wl_1_33 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2038 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_9 wl_1_9
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1326 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_17
+ wl_1_17 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2027 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_20 wl_1_20
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1315 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_28
+ wl_1_28 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2016 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_31 wl_1_31
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1304 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_39
+ wl_1_39 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2005 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_42 wl_1_42
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1348 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_59
+ wl_1_59 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1337 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_6
+ wl_1_6 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1359 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_48
+ wl_1_48 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_7 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_56
+ wl_1_56 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_712 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_55
+ wl_1_55 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_701 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_2
+ wl_1_2 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_756 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_11
+ wl_1_11 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_745 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_22
+ wl_1_22 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_734 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_33
+ wl_1_33 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_723 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_44
+ wl_1_44 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1860 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_59 wl_1_59
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_778 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_53
+ wl_1_53 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_767 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_0
+ wl_1_0 vdd_uq382 sky130_fd_bd_sram__openram_dp_cell_767/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_767/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1882 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_37 wl_1_37
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_789 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_42
+ wl_1_42 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1871 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_48 wl_1_48
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1893 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_26 wl_1_26
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_68 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_59
+ wl_1_59 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1156 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_59
+ wl_1_59 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_13 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_50
+ wl_1_50 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1101 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_50
+ wl_1_50 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_79 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_48
+ wl_1_48 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_57 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_6
+ wl_1_6 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1145 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_6
+ wl_1_6 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1134 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_17
+ wl_1_17 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_46 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_17
+ wl_1_17 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1123 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_28
+ wl_1_28 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_35 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_28
+ wl_1_28 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1112 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_39
+ wl_1_39 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_24 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_39
+ wl_1_39 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1167 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_48
+ wl_1_48 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1189 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_26
+ wl_1_26 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1178 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_37
+ wl_1_37 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_520 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_55
+ wl_1_55 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_586 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_53
+ wl_1_53 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_575 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_0
+ wl_1_0 vdd_uq286 sky130_fd_bd_sram__openram_dp_cell_575/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_575/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_564 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_11
+ wl_1_11 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_553 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_22
+ wl_1_22 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_542 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_33
+ wl_1_33 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_597 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_42
+ wl_1_42 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_531 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_44
+ wl_1_44 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1690 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_37 wl_1_37
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_394 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_53
+ wl_1_53 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_383 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_0
+ wl_1_0 vdd_uq190 sky130_fd_bd_sram__openram_dp_cell_383/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_383/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_372 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_11
+ wl_1_11 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_361 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_22
+ wl_1_22 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_350 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_33
+ wl_1_33 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_191 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_0
+ wl_1_0 vdd_uq94 sky130_fd_bd_sram__openram_dp_cell_191/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_191/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_180 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_11
+ wl_1_11 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1508 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_27 wl_1_27
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1519 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_16 wl_1_16
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_905 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_54
+ wl_1_54 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_949 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_10
+ wl_1_10 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_938 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_21
+ wl_1_21 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_927 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_32
+ wl_1_32 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_916 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_43
+ wl_1_43 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1349 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_58
+ wl_1_58 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2039 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_8 wl_1_8
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1338 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_5
+ wl_1_5 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1327 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_16
+ wl_1_16 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2028 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_19 wl_1_19
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1316 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_27
+ wl_1_27 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2017 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_30 wl_1_30
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1305 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_38
+ wl_1_38 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2006 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_41 wl_1_41
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_8 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_55
+ wl_1_55 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_768 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_63
+ wl_1_63 vdd_uq414 sky130_fd_bd_sram__openram_dp_cell_768/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_768/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_713 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_54
+ wl_1_54 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_779 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_52
+ wl_1_52 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_757 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_10
+ wl_1_10 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_702 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_1
+ wl_1_1 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_746 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_21
+ wl_1_21 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_735 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_32
+ wl_1_32 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_724 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_43
+ wl_1_43 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1861 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_58 wl_1_58
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1850 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_5 wl_1_5
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1894 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_25 wl_1_25
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1883 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_36 wl_1_36
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1872 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_47 wl_1_47
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_14 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_49
+ wl_1_49 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_69 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_58
+ wl_1_58 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1157 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_58
+ wl_1_58 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1102 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_49
+ wl_1_49 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_58 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_5
+ wl_1_5 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1146 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_5
+ wl_1_5 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1135 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_16
+ wl_1_16 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_47 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_16
+ wl_1_16 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1124 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_27
+ wl_1_27 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_36 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_27
+ wl_1_27 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1179 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_36
+ wl_1_36 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1113 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_38
+ wl_1_38 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_25 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_38
+ wl_1_38 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1168 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_47
+ wl_1_47 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_576 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_63
+ wl_1_63 vdd_uq318 sky130_fd_bd_sram__openram_dp_cell_576/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_576/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_521 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_54
+ wl_1_54 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_587 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_52
+ wl_1_52 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_565 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_10
+ wl_1_10 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_510 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_1
+ wl_1_1 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_554 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_21
+ wl_1_21 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_543 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_32
+ wl_1_32 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_598 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_41
+ wl_1_41 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_532 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_43
+ wl_1_43 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1691 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_36 wl_1_36
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1680 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_47 wl_1_47
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_340 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_43
+ wl_1_43 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_384 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_63
+ wl_1_63 vdd_uq222 sky130_fd_bd_sram__openram_dp_cell_384/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_384/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_395 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_52
+ wl_1_52 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_373 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_10
+ wl_1_10 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_362 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_21
+ wl_1_21 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_351 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_32
+ wl_1_32 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_181 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_10
+ wl_1_10 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_170 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_21
+ wl_1_21 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_192 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_63
+ wl_1_63 vdd_uq99 sky130_fd_bd_sram__openram_dp_cell_192/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_192/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1509 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_26 wl_1_26
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_906 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_53
+ wl_1_53 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_939 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_20
+ wl_1_20 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_928 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_31
+ wl_1_31 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_917 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_42
+ wl_1_42 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1339 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_4
+ wl_1_4 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1328 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_15
+ wl_1_15 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2029 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_18 wl_1_18
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1317 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_26
+ wl_1_26 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2018 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_29 wl_1_29
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1306 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_37
+ wl_1_37 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2007 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_40 wl_1_40
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_9 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_54
+ wl_1_54 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_769 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_62
+ wl_1_62 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_714 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_53
+ wl_1_53 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_758 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_9
+ wl_1_9 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_703 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_0
+ wl_1_0 vdd_uq350 sky130_fd_bd_sram__openram_dp_cell_703/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_703/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_747 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_20
+ wl_1_20 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_736 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_31
+ wl_1_31 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_725 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_42
+ wl_1_42 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1862 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_57 wl_1_57
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1851 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_4 wl_1_4
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1840 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_15 wl_1_15
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1895 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_24 wl_1_24
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1884 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_35 wl_1_35
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1873 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_46 wl_1_46
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_15 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_48
+ wl_1_48 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_48 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_15
+ wl_1_15 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_37 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_26
+ wl_1_26 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_26 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_37
+ wl_1_37 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1158 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_57
+ wl_1_57 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_59 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_4
+ wl_1_4 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1147 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_4
+ wl_1_4 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1136 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_15
+ wl_1_15 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1125 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_26
+ wl_1_26 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1114 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_37
+ wl_1_37 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1169 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_46
+ wl_1_46 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1103 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_48
+ wl_1_48 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_522 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_53
+ wl_1_53 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_511 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_0
+ wl_1_0 vdd_uq254 sky130_fd_bd_sram__openram_dp_cell_511/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_511/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_500 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_11
+ wl_1_11 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_577 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_62
+ wl_1_62 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_588 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_51
+ wl_1_51 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_566 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_9
+ wl_1_9 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_555 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_20
+ wl_1_20 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_544 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_31
+ wl_1_31 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_599 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_40
+ wl_1_40 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_533 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_42
+ wl_1_42 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1670 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_57 wl_1_57
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1692 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_35 wl_1_35
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1681 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_46 wl_1_46
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_330 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_53
+ wl_1_53 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_374 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_9
+ wl_1_9 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_363 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_20
+ wl_1_20 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_352 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_31
+ wl_1_31 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_341 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_42
+ wl_1_42 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_385 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_62
+ wl_1_62 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_396 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_51
+ wl_1_51 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_193 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_62
+ wl_1_62 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_182 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_9
+ wl_1_9 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_171 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_20
+ wl_1_20 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_160 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_31
+ wl_1_31 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_907 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_52
+ wl_1_52 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_929 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_30
+ wl_1_30 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_918 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_41
+ wl_1_41 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2019 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_28 wl_1_28
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2008 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_39 wl_1_39
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1329 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_14
+ wl_1_14 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1318 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_25
+ wl_1_25 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1307 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_36
+ wl_1_36 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_704 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_63
+ wl_1_63 vdd_uq382 sky130_fd_bd_sram__openram_dp_cell_704/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_704/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_715 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_52
+ wl_1_52 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_759 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_8
+ wl_1_8 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_748 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_19
+ wl_1_19 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1830 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_25 wl_1_25
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_737 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_30
+ wl_1_30 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_726 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_41
+ wl_1_41 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1863 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_56 wl_1_56
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1852 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_3 wl_1_3
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1841 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_14 wl_1_14
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1896 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_23 wl_1_23
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1885 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_34 wl_1_34
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1874 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_45 wl_1_45
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_16 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_47
+ wl_1_47 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_49 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_14
+ wl_1_14 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_38 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_25
+ wl_1_25 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1115 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_36
+ wl_1_36 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_27 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_36
+ wl_1_36 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1104 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_47
+ wl_1_47 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1159 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_56
+ wl_1_56 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1148 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_3
+ wl_1_3 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1137 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_14
+ wl_1_14 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1126 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_25
+ wl_1_25 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_512 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_63
+ wl_1_63 vdd_uq286 sky130_fd_bd_sram__openram_dp_cell_512/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_512/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_523 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_52
+ wl_1_52 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_501 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_10
+ wl_1_10 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_556 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_19
+ wl_1_19 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_545 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_30
+ wl_1_30 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_534 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_41
+ wl_1_41 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_578 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_61
+ wl_1_61 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1671 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_56 wl_1_56
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_589 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_50
+ wl_1_50 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_567 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_8
+ wl_1_8 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1660 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_3 wl_1_3
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1693 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_34 wl_1_34
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1682 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_45 wl_1_45
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_320 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_63
+ wl_1_63 vdd_uq190 sky130_fd_bd_sram__openram_dp_cell_320/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_320/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_386 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_61
+ wl_1_61 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_331 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_52
+ wl_1_52 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_397 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_50
+ wl_1_50 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_375 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_8
+ wl_1_8 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_364 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_19
+ wl_1_19 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_353 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_30
+ wl_1_30 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_342 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_41
+ wl_1_41 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1490 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_45 wl_1_45
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_194 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_61
+ wl_1_61 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_183 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_8
+ wl_1_8 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_172 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_19
+ wl_1_19 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_161 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_30
+ wl_1_30 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_150 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_41
+ wl_1_41 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_908 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_51
+ wl_1_51 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_919 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_40
+ wl_1_40 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1308 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_35
+ wl_1_35 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_2009 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_38 wl_1_38
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1319 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_24
+ wl_1_24 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_705 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_62
+ wl_1_62 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_716 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_51
+ wl_1_51 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_738 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_29
+ wl_1_29 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_727 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_40
+ wl_1_40 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1853 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_2 wl_1_2
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1842 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_13 wl_1_13
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_749 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_18
+ wl_1_18 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1831 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_24 wl_1_24
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1820 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_35 wl_1_35
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1864 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_55 wl_1_55
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1897 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_22 wl_1_22
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1886 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_33 wl_1_33
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1875 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_44 wl_1_44
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1149 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_2
+ wl_1_2 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1138 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_13
+ wl_1_13 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1127 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_24
+ wl_1_24 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_39 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_24
+ wl_1_24 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1116 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_35
+ wl_1_35 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_28 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_35
+ wl_1_35 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1105 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_46
+ wl_1_46 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_17 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_46
+ wl_1_46 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_513 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_62
+ wl_1_62 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_579 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_60
+ wl_1_60 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_524 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_51
+ wl_1_51 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_502 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_9
+ wl_1_9 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_568 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_7
+ wl_1_7 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_557 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_18
+ wl_1_18 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_546 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_29
+ wl_1_29 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_535 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_40
+ wl_1_40 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1672 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_55 wl_1_55
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1661 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_2 wl_1_2
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1650 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_13 wl_1_13
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1694 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_33 wl_1_33
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1683 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_44 wl_1_44
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_321 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_62
+ wl_1_62 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_387 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_60
+ wl_1_60 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_332 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_51
+ wl_1_51 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_398 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_49
+ wl_1_49 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_310 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_9
+ wl_1_9 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_376 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_7
+ wl_1_7 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_365 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_18
+ wl_1_18 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_354 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_29
+ wl_1_29 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_343 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_40
+ wl_1_40 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1480 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_55 wl_1_55
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1491 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_44 wl_1_44
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_140 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_51
+ wl_1_51 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_195 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_60
+ wl_1_60 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_184 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_7
+ wl_1_7 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_173 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_18
+ wl_1_18 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_162 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_29
+ wl_1_29 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_151 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_40
+ wl_1_40 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_909 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_50
+ wl_1_50 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1309 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_34
+ wl_1_34 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_706 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_61
+ wl_1_61 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_717 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_50
+ wl_1_50 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_739 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_28
+ wl_1_28 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_728 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_39
+ wl_1_39 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1865 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_54 wl_1_54
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1843 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_12 wl_1_12
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1854 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_1 wl_1_1
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1832 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_23 wl_1_23
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1887 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_32 wl_1_32
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1821 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_34 wl_1_34
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1876 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_43 wl_1_43
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1810 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_45 wl_1_45
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1898 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_21 wl_1_21
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1139 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_12
+ wl_1_12 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1128 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_23
+ wl_1_23 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1117 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_34
+ wl_1_34 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_29 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_34
+ wl_1_34 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1106 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_45
+ wl_1_45 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_18 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_45
+ wl_1_45 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_514 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_61
+ wl_1_61 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_525 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_50
+ wl_1_50 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_503 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_8
+ wl_1_8 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_569 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_6
+ wl_1_6 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_558 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_17
+ wl_1_17 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_547 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_28
+ wl_1_28 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_536 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_39
+ wl_1_39 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1673 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_54 wl_1_54
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1651 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_12 wl_1_12
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1662 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_1 wl_1_1
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1640 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_23 wl_1_23
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1695 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_32 wl_1_32
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1684 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_43 wl_1_43
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_322 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_61
+ wl_1_61 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_311 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_8
+ wl_1_8 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_300 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_19
+ wl_1_19 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_388 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_59
+ wl_1_59 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_333 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_50
+ wl_1_50 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_399 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_48
+ wl_1_48 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_377 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_6
+ wl_1_6 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_366 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_17
+ wl_1_17 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_355 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_28
+ wl_1_28 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_344 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_39
+ wl_1_39 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1481 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_54 wl_1_54
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1470 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_1 wl_1_1
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1492 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_43 wl_1_43
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_130 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_61
+ wl_1_61 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_141 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_50
+ wl_1_50 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_163 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_28
+ wl_1_28 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_152 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_39
+ wl_1_39 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_196 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_59
+ wl_1_59 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_185 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_6
+ wl_1_6 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_174 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_17
+ wl_1_17 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_707 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_60
+ wl_1_60 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_718 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_49
+ wl_1_49 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_729 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_38
+ wl_1_38 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1800 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_55 wl_1_55
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1866 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_53 wl_1_53
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1844 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_11 wl_1_11
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1855 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_0 wl_1_0
+ vdd_uq926 sky130_fd_bd_sram__openram_dp_cell_1855/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1855/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1899 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_20 wl_1_20
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1833 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_22 wl_1_22
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1888 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_31 wl_1_31
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1822 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_33 wl_1_33
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1877 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_42 wl_1_42
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1811 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_44 wl_1_44
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_19 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_44
+ wl_1_44 vdd bl_1_31 br_1_31 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1129 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_22
+ wl_1_22 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1118 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_33
+ wl_1_33 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1107 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_44
+ wl_1_44 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_504 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_7
+ wl_1_7 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_515 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_60
+ wl_1_60 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_526 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_49
+ wl_1_49 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_559 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_16
+ wl_1_16 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_548 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_27
+ wl_1_27 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_537 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_38
+ wl_1_38 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1674 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_53 wl_1_53
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1652 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_11 wl_1_11
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1663 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_0 wl_1_0
+ vdd_uq830 sky130_fd_bd_sram__openram_dp_cell_1663/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1663/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1641 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_22 wl_1_22
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1696 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_31 wl_1_31
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1630 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_33 wl_1_33
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1685 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_42 wl_1_42
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_323 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_60
+ wl_1_60 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_334 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_49
+ wl_1_49 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_312 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_7
+ wl_1_7 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_301 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_18
+ wl_1_18 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_356 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_27
+ wl_1_27 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_345 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_38
+ wl_1_38 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_389 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_58
+ wl_1_58 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1460 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_11 wl_1_11
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_378 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_5
+ wl_1_5 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1471 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_0 wl_1_0
+ vdd_uq734 sky130_fd_bd_sram__openram_dp_cell_1471/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1471/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_367 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_16
+ wl_1_16 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1482 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_53 wl_1_53
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1493 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_42 wl_1_42
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_890 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_5
+ wl_1_5 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_131 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_60
+ wl_1_60 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_197 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_58
+ wl_1_58 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_142 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_49
+ wl_1_49 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_120 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_7
+ wl_1_7 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_186 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_5
+ wl_1_5 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_175 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_16
+ wl_1_16 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_164 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_27
+ wl_1_27 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_153 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_38
+ wl_1_38 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1290 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_53
+ wl_1_53 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_708 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_59
+ wl_1_59 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1801 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_54 wl_1_54
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_719 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_48
+ wl_1_48 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1812 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_43 wl_1_43
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1856 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_63 wl_1_63
+ vdd_uq958 sky130_fd_bd_sram__openram_dp_cell_1856/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1856/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1867 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_52 wl_1_52
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1845 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_10 wl_1_10
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1834 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_21 wl_1_21
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1889 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_30 wl_1_30
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1823 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_32 wl_1_32
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1878 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_41 wl_1_41
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1119 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_32
+ wl_1_32 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1108 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_43
+ wl_1_43 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_516 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_59
+ wl_1_59 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_527 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_48
+ wl_1_48 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_505 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_6
+ wl_1_6 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_538 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_37
+ wl_1_37 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1653 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_10 wl_1_10
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1642 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_21 wl_1_21
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_549 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_26
+ wl_1_26 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1631 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_32 wl_1_32
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1620 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_43 wl_1_43
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1664 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_63 wl_1_63
+ vdd_uq862 sky130_fd_bd_sram__openram_dp_cell_1664/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1664/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1675 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_52 wl_1_52
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1697 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_30 wl_1_30
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1686 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_41 wl_1_41
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_324 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_59
+ wl_1_59 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_335 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_48
+ wl_1_48 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_313 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_6
+ wl_1_6 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_379 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_4
+ wl_1_4 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_368 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_15
+ wl_1_15 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_302 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_17
+ wl_1_17 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_357 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_26
+ wl_1_26 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_346 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_37
+ wl_1_37 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1472 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_63 wl_1_63
+ vdd_uq766 sky130_fd_bd_sram__openram_dp_cell_1472/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1472/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1483 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_52 wl_1_52
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1461 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_10 wl_1_10
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1450 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_21 wl_1_21
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1494 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_41 wl_1_41
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_891 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_4
+ wl_1_4 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_880 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_15
+ wl_1_15 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_132 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_59
+ wl_1_59 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_198 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_57
+ wl_1_57 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_143 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_48
+ wl_1_48 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_121 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_6
+ wl_1_6 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_187 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_4
+ wl_1_4 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_176 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_15
+ wl_1_15 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_110 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_17
+ wl_1_17 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_165 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_26
+ wl_1_26 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_154 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_37
+ wl_1_37 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1280 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_63
+ wl_1_63 vdd_uq670 sky130_fd_bd_sram__openram_dp_cell_1280/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1280/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1291 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_52
+ wl_1_52 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_709 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_58
+ wl_1_58 vdd_uq382 bl_1_20 br_1_20 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1802 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_53 wl_1_53
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1835 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_20 wl_1_20
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1824 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_31 wl_1_31
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1813 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_42 wl_1_42
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1857 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_62 wl_1_62
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1868 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_51 wl_1_51
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1846 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_9 wl_1_9
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1879 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_40 wl_1_40
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1109 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_42
+ wl_1_42 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_517 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_58
+ wl_1_58 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_528 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_47
+ wl_1_47 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_506 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_5
+ wl_1_5 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_539 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_36
+ wl_1_36 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1665 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_62 wl_1_62
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1610 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_53 wl_1_53
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1676 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_51 wl_1_51
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1654 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_9 wl_1_9
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1643 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_20 wl_1_20
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1632 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_31 wl_1_31
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1687 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_40 wl_1_40
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1621 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_42 wl_1_42
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1698 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_29 wl_1_29
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_325 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_58
+ wl_1_58 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_336 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_47
+ wl_1_47 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_314 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_5
+ wl_1_5 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_369 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_14
+ wl_1_14 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_303 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_16
+ wl_1_16 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_358 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_25
+ wl_1_25 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_347 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_36
+ wl_1_36 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1473 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_62 wl_1_62
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1484 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_51 wl_1_51
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1462 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_9 wl_1_9
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1451 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_20 wl_1_20
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1440 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_31 wl_1_31
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1495 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_40 wl_1_40
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_892 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_3
+ wl_1_3 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_881 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_14
+ wl_1_14 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_870 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_25
+ wl_1_25 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_122 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_5
+ wl_1_5 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_111 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_16
+ wl_1_16 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_100 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_27
+ wl_1_27 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_133 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_58
+ wl_1_58 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_199 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_56
+ wl_1_56 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_144 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_47
+ wl_1_47 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_188 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_3
+ wl_1_3 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_177 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_14
+ wl_1_14 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_166 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_25
+ wl_1_25 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_155 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_36
+ wl_1_36 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1281 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_62
+ wl_1_62 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1292 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_51
+ wl_1_51 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1270 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_9
+ wl_1_9 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1858 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_61 wl_1_61
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1803 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_52 wl_1_52
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1869 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_50 wl_1_50
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1847 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_8 wl_1_8
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1836 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_19 wl_1_19
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1825 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_30 wl_1_30
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1814 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_41 wl_1_41
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_518 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_57
+ wl_1_57 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_507 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_4
+ wl_1_4 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_529 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_46
+ wl_1_46 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1600 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_63 wl_1_63
+ vdd_uq830 sky130_fd_bd_sram__openram_dp_cell_1600/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1600/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1666 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_61 wl_1_61
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1611 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_52 wl_1_52
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1677 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_50 wl_1_50
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1655 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_8 wl_1_8
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1644 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_19 wl_1_19
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1699 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_28 wl_1_28
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1633 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_30 wl_1_30
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1688 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_39 wl_1_39
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1622 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_41 wl_1_41
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_304 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_15
+ wl_1_15 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_326 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_57
+ wl_1_57 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_315 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_4
+ wl_1_4 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_359 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_24
+ wl_1_24 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_348 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_35
+ wl_1_35 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_337 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_46
+ wl_1_46 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1474 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_61 wl_1_61
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1485 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_50 wl_1_50
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1463 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_8 wl_1_8
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1452 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_19 wl_1_19
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1441 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_30 wl_1_30
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1496 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_39 wl_1_39
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1430 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_41 wl_1_41
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_860 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_35
+ wl_1_35 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_893 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_2
+ wl_1_2 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_882 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_13
+ wl_1_13 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_871 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_24
+ wl_1_24 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_134 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_57
+ wl_1_57 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_123 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_4
+ wl_1_4 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_112 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_15
+ wl_1_15 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_101 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_26
+ wl_1_26 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_145 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_46
+ wl_1_46 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1271 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_8
+ wl_1_8 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_189 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_2
+ wl_1_2 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_178 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_13
+ wl_1_13 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1260 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_19
+ wl_1_19 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_167 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_24
+ wl_1_24 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_156 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_35
+ wl_1_35 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1282 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_61
+ wl_1_61 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1293 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_50
+ wl_1_50 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_690 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_13
+ wl_1_13 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1090 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_61
+ wl_1_61 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1859 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_60 wl_1_60
+ vdd_uq958 bl_1_2 br_1_2 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1804 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_51 wl_1_51
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1848 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_7 wl_1_7
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1837 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_18 wl_1_18
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1826 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_29 wl_1_29
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1815 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_40 wl_1_40
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1601 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_62 wl_1_62
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_519 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_56
+ wl_1_56 vdd_uq286 bl_1_23 br_1_23 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_508 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_3
+ wl_1_3 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1667 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_60 wl_1_60
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1612 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_51 wl_1_51
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1678 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_49 wl_1_49
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1656 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_7 wl_1_7
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1645 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_18 wl_1_18
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1634 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_29 wl_1_29
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1689 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_38 wl_1_38
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1623 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_40 wl_1_40
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_327 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_56
+ wl_1_56 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_316 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_3
+ wl_1_3 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_305 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_14
+ wl_1_14 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_338 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_45
+ wl_1_45 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1420 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_51 wl_1_51
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1453 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_18 wl_1_18
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1442 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_29 wl_1_29
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_349 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_34
+ wl_1_34 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1431 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_40 wl_1_40
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1475 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_60 wl_1_60
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1486 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_49 wl_1_49
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1464 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_7 wl_1_7
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1497 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_38 wl_1_38
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_894 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_1
+ wl_1_1 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_883 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_12
+ wl_1_12 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_872 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_23
+ wl_1_23 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_861 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_34
+ wl_1_34 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_850 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_45
+ wl_1_45 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_135 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_56
+ wl_1_56 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_124 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_3
+ wl_1_3 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_179 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_12
+ wl_1_12 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_113 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_14
+ wl_1_14 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_168 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_23
+ wl_1_23 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_102 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_25
+ wl_1_25 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_157 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_34
+ wl_1_34 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_146 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_45
+ wl_1_45 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1283 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_60
+ wl_1_60 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1294 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_49
+ wl_1_49 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1272 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_7
+ wl_1_7 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1261 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_18
+ wl_1_18 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1250 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_29
+ wl_1_29 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_691 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_12
+ wl_1_12 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_680 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_23
+ wl_1_23 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1091 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_60
+ wl_1_60 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1080 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_7
+ wl_1_7 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1805 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_50 wl_1_50
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1849 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_6 wl_1_6
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1838 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_17 wl_1_17
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1827 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_28 wl_1_28
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1816 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_39 wl_1_39
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_509 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_2
+ wl_1_2 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1602 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_61 wl_1_61
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1613 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_50 wl_1_50
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1635 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_28 wl_1_28
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1624 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_39 wl_1_39
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1668 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_59 wl_1_59
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1657 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_6 wl_1_6
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1646 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_17 wl_1_17
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1679 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_48 wl_1_48
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_328 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_55
+ wl_1_55 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_317 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_2
+ wl_1_2 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_306 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_13
+ wl_1_13 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_339 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_44
+ wl_1_44 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1410 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_61 wl_1_61
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1476 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_59 wl_1_59
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1421 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_50 wl_1_50
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1465 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_6 wl_1_6
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1454 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_17 wl_1_17
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1443 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_28 wl_1_28
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1432 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_39 wl_1_39
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1487 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_48 wl_1_48
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1498 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_37 wl_1_37
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_840 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_55
+ wl_1_55 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_895 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_0
+ wl_1_0 vdd_uq446 sky130_fd_bd_sram__openram_dp_cell_895/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_895/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_884 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_11
+ wl_1_11 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_873 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_22
+ wl_1_22 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_862 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_33
+ wl_1_33 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_851 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_44
+ wl_1_44 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_136 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_55
+ wl_1_55 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_125 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_2
+ wl_1_2 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_114 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_13
+ wl_1_13 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_169 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_22
+ wl_1_22 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_103 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_24
+ wl_1_24 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_158 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_33
+ wl_1_33 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_147 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_44
+ wl_1_44 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1284 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_59
+ wl_1_59 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1273 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_6
+ wl_1_6 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1262 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_17
+ wl_1_17 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1251 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_28
+ wl_1_28 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1240 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_39
+ wl_1_39 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1295 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_48
+ wl_1_48 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_692 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_11
+ wl_1_11 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_681 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_22
+ wl_1_22 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_670 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_33
+ wl_1_33 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1092 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_59
+ wl_1_59 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1081 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_6
+ wl_1_6 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1070 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_17
+ wl_1_17 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1806 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_49 wl_1_49
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1817 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_38 wl_1_38
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1839 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_16 wl_1_16
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1828 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_27 wl_1_27
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1603 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_60 wl_1_60
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1669 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_58 wl_1_58
+ vdd_uq862 bl_1_5 br_1_5 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1614 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_49 wl_1_49
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1658 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_5 wl_1_5
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1647 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_16 wl_1_16
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1636 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_27 wl_1_27
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1625 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_38 wl_1_38
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_329 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_54
+ wl_1_54 vdd_uq190 bl_1_26 br_1_26 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_318 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_1
+ wl_1_1 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_307 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_12
+ wl_1_12 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1411 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_60 wl_1_60
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1477 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_58 wl_1_58
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1422 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_49 wl_1_49
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1400 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_7
+ wl_1_7 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1466 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_5 wl_1_5
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1455 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_16 wl_1_16
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1444 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_27 wl_1_27
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1499 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_36 wl_1_36
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1433 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_38 wl_1_38
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1488 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_47 wl_1_47
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_896 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_63
+ wl_1_63 vdd_uq478 sky130_fd_bd_sram__openram_dp_cell_896/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_896/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_841 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_54
+ wl_1_54 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_885 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_10
+ wl_1_10 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_830 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_1
+ wl_1_1 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_874 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_21
+ wl_1_21 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_863 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_32
+ wl_1_32 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_852 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_43
+ wl_1_43 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_104 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_23
+ wl_1_23 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_137 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_54
+ wl_1_54 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_126 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_1
+ wl_1_1 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_115 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_12
+ wl_1_12 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_159 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_32
+ wl_1_32 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_148 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_43
+ wl_1_43 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1285 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_58
+ wl_1_58 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1230 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_49
+ wl_1_49 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1274 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_5
+ wl_1_5 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1263 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_16
+ wl_1_16 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1252 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_27
+ wl_1_27 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1241 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_38
+ wl_1_38 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1296 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_47
+ wl_1_47 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_693 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_10
+ wl_1_10 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_682 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_21
+ wl_1_21 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_671 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_32
+ wl_1_32 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_660 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_43
+ wl_1_43 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1060 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_27
+ wl_1_27 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1093 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_58
+ wl_1_58 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1082 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_5
+ wl_1_5 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1071 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_16
+ wl_1_16 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_490 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_21
+ wl_1_21 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1829 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_26 wl_1_26
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1818 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_37 wl_1_37
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1807 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_48 wl_1_48
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1604 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_59 wl_1_59
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1659 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_4 wl_1_4
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1648 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_15 wl_1_15
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1637 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_26 wl_1_26
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1626 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_37 wl_1_37
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1615 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_48 wl_1_48
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1401 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_6
+ wl_1_6 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_319 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_0
+ wl_1_0 vdd_uq158 sky130_fd_bd_sram__openram_dp_cell_319/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_319/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_308 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_11
+ wl_1_11 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1412 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_59 wl_1_59
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1478 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_57 wl_1_57
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1467 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_4 wl_1_4
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1456 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_15 wl_1_15
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1445 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_26 wl_1_26
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1434 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_37 wl_1_37
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1489 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_46 wl_1_46
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1423 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_48 wl_1_48
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_842 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_53
+ wl_1_53 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_831 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_0
+ wl_1_0 vdd_uq414 sky130_fd_bd_sram__openram_dp_cell_831/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_831/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_820 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_11
+ wl_1_11 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_897 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_62
+ wl_1_62 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_886 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_9
+ wl_1_9 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_875 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_20
+ wl_1_20 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_864 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_31
+ wl_1_31 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_853 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_42
+ wl_1_42 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1990 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_57 wl_1_57
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_127 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_0
+ wl_1_0 vdd_uq62 sky130_fd_bd_sram__openram_dp_cell_127/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_127/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_116 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_11
+ wl_1_11 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_105 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_22
+ wl_1_22 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1220 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_59
+ wl_1_59 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_138 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_53
+ wl_1_53 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1253 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_26
+ wl_1_26 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1242 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_37
+ wl_1_37 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_149 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_42
+ wl_1_42 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1231 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_48
+ wl_1_48 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1286 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_57
+ wl_1_57 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1275 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_4
+ wl_1_4 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1264 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_15
+ wl_1_15 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1297 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_46
+ wl_1_46 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_650 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_53
+ wl_1_53 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_683 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_20
+ wl_1_20 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_672 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_31
+ wl_1_31 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_661 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_42
+ wl_1_42 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_694 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_9
+ wl_1_9 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1094 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_57
+ wl_1_57 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1083 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_4
+ wl_1_4 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1072 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_15
+ wl_1_15 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1061 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_26
+ wl_1_26 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1050 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_37
+ wl_1_37 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_491 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_20
+ wl_1_20 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_480 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_31
+ wl_1_31 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1819 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_36 wl_1_36
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1808 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_47 wl_1_47
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1605 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_58 wl_1_58
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1649 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_14 wl_1_14
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1638 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_25 wl_1_25
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1627 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_36 wl_1_36
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1616 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_47 wl_1_47
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_309 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_10
+ wl_1_10 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1413 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_58 wl_1_58
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1402 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_5
+ wl_1_5 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1435 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_36 wl_1_36
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1424 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_47 wl_1_47
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1479 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_56 wl_1_56
+ vdd_uq766 bl_1_8 br_1_8 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1468 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_3 wl_1_3
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1457 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_14 wl_1_14
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1446 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_25 wl_1_25
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_832 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_63
+ wl_1_63 vdd_uq446 sky130_fd_bd_sram__openram_dp_cell_832/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_832/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_843 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_52
+ wl_1_52 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_821 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_10
+ wl_1_10 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_810 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_21
+ wl_1_21 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_865 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_30
+ wl_1_30 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_854 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_41
+ wl_1_41 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_898 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_61
+ wl_1_61 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1991 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_56 wl_1_56
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_887 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_8
+ wl_1_8 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1980 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_3 wl_1_3
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_876 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_19
+ wl_1_19 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_128 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_63
+ wl_1_63 vdd_uq94 sky130_fd_bd_sram__openram_dp_cell_128/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_128/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_139 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_52
+ wl_1_52 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_117 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_10
+ wl_1_10 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_106 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_21
+ wl_1_21 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1221 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_58
+ wl_1_58 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1210 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_5
+ wl_1_5 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1276 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_3
+ wl_1_3 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1265 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_14
+ wl_1_14 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1254 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_25
+ wl_1_25 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1243 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_36
+ wl_1_36 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1232 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_47
+ wl_1_47 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1287 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_56
+ wl_1_56 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1298 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_45
+ wl_1_45 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_640 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_63
+ wl_1_63 vdd_uq350 sky130_fd_bd_sram__openram_dp_cell_640/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_640/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_651 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_52
+ wl_1_52 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_695 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_8
+ wl_1_8 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_684 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_19
+ wl_1_19 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_673 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_30
+ wl_1_30 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_662 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_41
+ wl_1_41 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1095 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_56
+ wl_1_56 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1084 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_3
+ wl_1_3 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1073 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_14
+ wl_1_14 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1062 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_25
+ wl_1_25 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1051 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_36
+ wl_1_36 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1040 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_47
+ wl_1_47 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_492 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_19
+ wl_1_19 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_481 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_30
+ wl_1_30 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_470 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_41
+ wl_1_41 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1809 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_46 wl_1_46
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1606 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_57 wl_1_57
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1617 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_46 wl_1_46
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1639 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_24 wl_1_24
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1628 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_35 wl_1_35
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1414 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_57 wl_1_57
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1403 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_4
+ wl_1_4 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1469 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_2 wl_1_2
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1458 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_13 wl_1_13
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1447 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_24 wl_1_24
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1436 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_35 wl_1_35
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1425 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_46 wl_1_46
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_833 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_62
+ wl_1_62 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_899 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_60
+ wl_1_60 vdd_uq478 bl_1_17 br_1_17 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_844 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_51
+ wl_1_51 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_822 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_9
+ wl_1_9 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_888 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_7
+ wl_1_7 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_877 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_18
+ wl_1_18 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_811 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_20
+ wl_1_20 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_866 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_29
+ wl_1_29 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_800 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_31
+ wl_1_31 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_855 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_40
+ wl_1_40 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1992 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_55 wl_1_55
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1981 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_2 wl_1_2
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1970 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_13 wl_1_13
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_129 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_62
+ wl_1_62 vdd_uq94 bl_1_29 br_1_29 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_118 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_9
+ wl_1_9 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_107 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_20
+ wl_1_20 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1222 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_57
+ wl_1_57 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1288 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_55
+ wl_1_55 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1211 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_4
+ wl_1_4 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1277 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_2
+ wl_1_2 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1266 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_13
+ wl_1_13 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1200 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_15
+ wl_1_15 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1255 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_24
+ wl_1_24 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1244 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_35
+ wl_1_35 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1299 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_44
+ wl_1_44 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1233 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_46
+ wl_1_46 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_641 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_62
+ wl_1_62 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_652 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_51
+ wl_1_51 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_630 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_9
+ wl_1_9 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_696 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_7
+ wl_1_7 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_685 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_18
+ wl_1_18 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_674 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_29
+ wl_1_29 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_663 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_40
+ wl_1_40 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1030 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_57
+ wl_1_57 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1096 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_55
+ wl_1_55 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1085 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_2
+ wl_1_2 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1074 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_13
+ wl_1_13 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1063 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_24
+ wl_1_24 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1052 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_35
+ wl_1_35 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1041 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_46
+ wl_1_46 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_460 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_51
+ wl_1_51 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_493 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_18
+ wl_1_18 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_482 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_29
+ wl_1_29 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_471 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_40
+ wl_1_40 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_290 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_29
+ wl_1_29 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1607 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_56 wl_1_56
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1629 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_34 wl_1_34
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1618 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_45 wl_1_45
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1415 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_56 wl_1_56
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1459 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_12 wl_1_12
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1404 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_3
+ wl_1_3 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1448 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_23 wl_1_23
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1437 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_34 wl_1_34
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1426 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_45 wl_1_45
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_834 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_61
+ wl_1_61 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_845 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_50
+ wl_1_50 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_823 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_8
+ wl_1_8 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_889 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_6
+ wl_1_6 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_878 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_17
+ wl_1_17 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_812 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_19
+ wl_1_19 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_867 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_28
+ wl_1_28 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_801 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_30
+ wl_1_30 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_856 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_39
+ wl_1_39 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1993 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_54 wl_1_54
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1971 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_12 wl_1_12
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1982 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_1 wl_1_1
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1960 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_23 wl_1_23
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_119 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_8
+ wl_1_8 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1201 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_14
+ wl_1_14 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_108 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_19
+ wl_1_19 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1223 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_56
+ wl_1_56 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1289 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_54
+ wl_1_54 vdd_uq670 bl_1_11 br_1_11 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1267 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_12
+ wl_1_12 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1212 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_3
+ wl_1_3 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1278 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_1
+ wl_1_1 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1256 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_23
+ wl_1_23 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1245 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_34
+ wl_1_34 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1234 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_45
+ wl_1_45 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_631 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_8
+ wl_1_8 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_620 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_19
+ wl_1_19 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_642 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_61
+ wl_1_61 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_653 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_50
+ wl_1_50 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_697 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_6
+ wl_1_6 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_686 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_17
+ wl_1_17 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_675 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_28
+ wl_1_28 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_664 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_39
+ wl_1_39 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1790 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_1 wl_1_1
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1031 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_56
+ wl_1_56 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1020 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_3
+ wl_1_3 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1042 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_45
+ wl_1_45 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1097 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_54
+ wl_1_54 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1075 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_12
+ wl_1_12 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1086 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_1
+ wl_1_1 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1064 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_23
+ wl_1_23 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1053 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_34
+ wl_1_34 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_450 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_61
+ wl_1_61 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_461 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_50
+ wl_1_50 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_483 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_28
+ wl_1_28 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_472 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_39
+ wl_1_39 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_494 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_17
+ wl_1_17 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_291 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_28
+ wl_1_28 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_280 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_39
+ wl_1_39 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1608 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_55 wl_1_55
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1619 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_44 wl_1_44
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1416 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_55 wl_1_55
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1405 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_2
+ wl_1_2 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1449 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_22 wl_1_22
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1438 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_33 wl_1_33
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1427 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_44 wl_1_44
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_824 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_7
+ wl_1_7 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_813 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_18
+ wl_1_18 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_802 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_29
+ wl_1_29 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_835 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_60
+ wl_1_60 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_846 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_49
+ wl_1_49 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_879 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_16
+ wl_1_16 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_868 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_27
+ wl_1_27 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_857 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_38
+ wl_1_38 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1994 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_53 wl_1_53
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1972 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_11 wl_1_11
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1983 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_0 wl_1_0
+ vdd_uq990 sky130_fd_bd_sram__openram_dp_cell_1983/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1983/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1961 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_22 wl_1_22
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1950 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_33 wl_1_33
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_109 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_18
+ wl_1_18 vdd_uq62 bl_1_30 br_1_30 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1224 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_55
+ wl_1_55 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1213 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_2
+ wl_1_2 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1202 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_13
+ wl_1_13 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1235 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_44
+ wl_1_44 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1268 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_11
+ wl_1_11 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1279 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_0
+ wl_1_0 vdd_uq638 sky130_fd_bd_sram__openram_dp_cell_1279/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1279/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1257 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_22
+ wl_1_22 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1246 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_33
+ wl_1_33 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_643 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_60
+ wl_1_60 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_654 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_49
+ wl_1_49 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_632 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_7
+ wl_1_7 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_621 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_18
+ wl_1_18 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_610 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_29
+ wl_1_29 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_665 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_38
+ wl_1_38 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1780 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_11 wl_1_11
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_698 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_5
+ wl_1_5 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_687 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_16
+ wl_1_16 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_676 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_27
+ wl_1_27 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1791 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_0 wl_1_0
+ vdd_uq894 sky130_fd_bd_sram__openram_dp_cell_1791/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1791/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1032 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_55
+ wl_1_55 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1076 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_11
+ wl_1_11 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1021 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_2
+ wl_1_2 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1010 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_13
+ wl_1_13 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1065 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_22
+ wl_1_22 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1054 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_33
+ wl_1_33 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1043 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_44
+ wl_1_44 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1098 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_53
+ wl_1_53 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1087 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_0
+ wl_1_0 vdd_uq542 sky130_fd_bd_sram__openram_dp_cell_1087/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1087/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_451 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_60
+ wl_1_60 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_462 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_49
+ wl_1_49 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_440 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_7
+ wl_1_7 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_495 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_16
+ wl_1_16 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_484 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_27
+ wl_1_27 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_473 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_38
+ wl_1_38 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_270 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_49
+ wl_1_49 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_292 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_27
+ wl_1_27 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_281 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_38
+ wl_1_38 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1609 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_54 wl_1_54
+ vdd_uq830 bl_1_6 br_1_6 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1417 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_54 wl_1_54
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1406 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_1
+ wl_1_1 vdd_uq702 bl_1_10 br_1_10 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1439 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_32 wl_1_32
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1428 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_43 wl_1_43
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_836 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_59
+ wl_1_59 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_847 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_48
+ wl_1_48 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_825 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_6
+ wl_1_6 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_814 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_17
+ wl_1_17 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_803 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_28
+ wl_1_28 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1973 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_10 wl_1_10
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1962 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_21 wl_1_21
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_869 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_26
+ wl_1_26 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1951 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_32 wl_1_32
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_858 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_37
+ wl_1_37 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1940 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_43 wl_1_43
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1984 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_63 wl_1_63
+ vdd_uq999 sky130_fd_bd_sram__openram_dp_cell_1984/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1984/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1995 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_52 wl_1_52
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1225 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_54
+ wl_1_54 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1203 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_12
+ wl_1_12 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1214 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_1
+ wl_1_1 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1258 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_21
+ wl_1_21 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1247 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_32
+ wl_1_32 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1236 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_43
+ wl_1_43 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1269 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_10
+ wl_1_10 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_644 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_59
+ wl_1_59 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_655 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_48
+ wl_1_48 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_633 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_6
+ wl_1_6 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_699 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_4
+ wl_1_4 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_688 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_15
+ wl_1_15 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_622 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_17
+ wl_1_17 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_677 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_26
+ wl_1_26 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_611 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_28
+ wl_1_28 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_666 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_37
+ wl_1_37 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_600 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_39
+ wl_1_39 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1792 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_63 wl_1_63
+ vdd_uq926 sky130_fd_bd_sram__openram_dp_cell_1792/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1792/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1781 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_10 wl_1_10
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1770 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_21 wl_1_21
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1088 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_63
+ wl_1_63 vdd_uq574 sky130_fd_bd_sram__openram_dp_cell_1088/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1088/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1033 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_54
+ wl_1_54 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1099 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_52
+ wl_1_52 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1077 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_10
+ wl_1_10 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1022 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_1
+ wl_1_1 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1011 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_12
+ wl_1_12 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1066 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_21
+ wl_1_21 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1000 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_23
+ wl_1_23 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1055 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_32
+ wl_1_32 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1044 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_43
+ wl_1_43 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_452 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_59
+ wl_1_59 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_463 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_48
+ wl_1_48 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_441 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_6
+ wl_1_6 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_496 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_15
+ wl_1_15 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_430 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_17
+ wl_1_17 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_485 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_26
+ wl_1_26 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_474 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_37
+ wl_1_37 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_260 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_59
+ wl_1_59 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_271 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_48
+ wl_1_48 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_293 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_26
+ wl_1_26 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_282 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_37
+ wl_1_37 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1418 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_53 wl_1_53
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1407 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_0
+ wl_1_0 vdd_uq702 sky130_fd_bd_sram__openram_dp_cell_1407/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1407/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1429 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_42 wl_1_42
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_837 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_58
+ wl_1_58 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_848 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_47
+ wl_1_47 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_826 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_5
+ wl_1_5 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_815 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_16
+ wl_1_16 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_804 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_27
+ wl_1_27 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_859 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_36
+ wl_1_36 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1985 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_62 wl_1_62
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1930 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_53 wl_1_53
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1996 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_51 wl_1_51
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1974 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_9 wl_1_9
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1963 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_20 wl_1_20
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1952 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_31 wl_1_31
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1941 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_42 wl_1_42
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1226 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_53
+ wl_1_53 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1204 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_11
+ wl_1_11 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1215 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_0
+ wl_1_0 vdd_uq606 sky130_fd_bd_sram__openram_dp_cell_1215/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1215/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1259 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_20
+ wl_1_20 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1248 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_31
+ wl_1_31 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1237 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_42
+ wl_1_42 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_645 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_58
+ wl_1_58 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_656 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_47
+ wl_1_47 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_634 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_5
+ wl_1_5 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_689 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_14
+ wl_1_14 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_623 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_16
+ wl_1_16 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_678 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_25
+ wl_1_25 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_612 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_27
+ wl_1_27 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_667 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_36
+ wl_1_36 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_601 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_38
+ wl_1_38 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1793 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_62 wl_1_62
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1782 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_9 wl_1_9
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1771 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_20 wl_1_20
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1760 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_31 wl_1_31
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1089 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_62
+ wl_1_62 vdd_uq574 bl_1_14 br_1_14 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1034 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_53
+ wl_1_53 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1078 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_9
+ wl_1_9 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1023 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_0
+ wl_1_0 vdd_uq510 sky130_fd_bd_sram__openram_dp_cell_1023/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1023/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1012 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_11
+ wl_1_11 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1067 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_20
+ wl_1_20 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1001 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_22
+ wl_1_22 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1056 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_31
+ wl_1_31 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1045 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_42
+ wl_1_42 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_431 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_16
+ wl_1_16 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_420 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_27
+ wl_1_27 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_453 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_58
+ wl_1_58 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_464 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_47
+ wl_1_47 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_442 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_5
+ wl_1_5 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_497 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_14
+ wl_1_14 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_486 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_25
+ wl_1_25 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_475 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_36
+ wl_1_36 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1590 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_9 wl_1_9
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_261 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_58
+ wl_1_58 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_272 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_47
+ wl_1_47 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_250 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_5
+ wl_1_5 vdd_uq99 bl_1_28 br_1_28 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_283 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_36
+ wl_1_36 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_294 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_25
+ wl_1_25 vdd_uq158 bl_1_27 br_1_27 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1408 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_63 wl_1_63
+ vdd_uq734 sky130_fd_bd_sram__openram_dp_cell_1408/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1408/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1419 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_52 wl_1_52
+ vdd_uq734 bl_1_9 br_1_9 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_838 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_57
+ wl_1_57 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_827 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_4
+ wl_1_4 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_816 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_15
+ wl_1_15 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_805 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_26
+ wl_1_26 vdd_uq414 bl_1_19 br_1_19 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_849 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_46
+ wl_1_46 vdd_uq446 bl_1_18 br_1_18 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1920 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_63 wl_1_63
+ vdd_uq990 sky130_fd_bd_sram__openram_dp_cell_1920/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1920/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1986 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_61 wl_1_61
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1931 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_52 wl_1_52
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1997 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_50 wl_1_50
+ vdd_uq999 bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1975 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_8 wl_1_8
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1964 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_19 wl_1_19
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1953 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_30 wl_1_30
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1942 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_41 wl_1_41
+ vdd_uq990 bl_1_1 br_1_1 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1216 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_63
+ wl_1_63 vdd_uq638 sky130_fd_bd_sram__openram_dp_cell_1216/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1216/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1227 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_52
+ wl_1_52 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1205 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_10
+ wl_1_10 vdd_uq606 bl_1_13 br_1_13 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1249 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_30
+ wl_1_30 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1238 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_41
+ wl_1_41 vdd_uq638 bl_1_12 br_1_12 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_613 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_26
+ wl_1_26 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_602 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_37
+ wl_1_37 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_646 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_57
+ wl_1_57 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_635 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_4
+ wl_1_4 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_624 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_15
+ wl_1_15 vdd_uq318 bl_1_22 br_1_22 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_679 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_24
+ wl_1_24 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_668 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_35
+ wl_1_35 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_657 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_46
+ wl_1_46 vdd_uq350 bl_1_21 br_1_21 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1794 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_61 wl_1_61
+ vdd_uq926 bl_1_3 br_1_3 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1783 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_8 wl_1_8
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1772 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_19 wl_1_19
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1761 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_30 wl_1_30
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1750 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_41 wl_1_41
+ vdd_uq894 bl_1_4 br_1_4 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1024 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_63
+ wl_1_63 vdd_uq542 sky130_fd_bd_sram__openram_dp_cell_1024/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_1024/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1013 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_10
+ wl_1_10 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1002 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_21
+ wl_1_21 vdd_uq510 bl_1_16 br_1_16 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1035 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_52
+ wl_1_52 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1079 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_8
+ wl_1_8 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1068 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_19
+ wl_1_19 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1057 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_30
+ wl_1_30 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1046 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_41
+ wl_1_41 vdd_uq542 bl_1_15 br_1_15 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_454 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_57
+ wl_1_57 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_443 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_4
+ wl_1_4 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_432 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_15
+ wl_1_15 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_421 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_26
+ wl_1_26 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_410 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_37
+ wl_1_37 vdd_uq222 bl_1_25 br_1_25 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_465 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_46
+ wl_1_46 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_498 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_13
+ wl_1_13 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1580 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_19 wl_1_19
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_487 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_24
+ wl_1_24 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_476 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_35
+ wl_1_35 vdd_uq254 bl_1_24 br_1_24 sky130_fd_bd_sram__openram_dp_cell
Xsky130_fd_bd_sram__openram_dp_cell_1591 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_8 wl_1_8
+ vdd_uq798 bl_1_7 br_1_7 sky130_fd_bd_sram__openram_dp_cell
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell_dummy gnd bl0 br0 bl1 br1 wl0 wl1 vdd a_38_n79#
+ w_144_n79# a_400_n79#
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=1.6583p pd=22.5u as=0.0504p ps=0.9u w=0.21u l=0.08u
X1 a_400_133# wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0504p ps=0.9u w=0.21u l=0.15u
X2 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X3 a_400_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.2768p ps=4u w=0.21u l=0.15u
X4 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X5 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X6 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.08u
X7 a_38_291# gnd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X8 br0 wl0 a_400_291# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0525p ps=0.92u w=0.21u l=0.15u
X9 gnd gnd a_400_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0525p ps=0.92u w=0.21u l=0.15u
X10 bl0 wl0 a_38_291# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0525p ps=0.92u w=0.21u l=0.15u
X11 gnd gnd a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0525p ps=0.92u w=0.21u l=0.15u
.ends

.subckt subbyte2_dummy_array br_1_0 bl_0_1 br_1_1 br_1_3 bl_0_4 bl_1_4 br_1_4 bl_1_5
+ br_0_5 br_1_5 bl_1_6 br_1_6 bl_0_7 bl_1_7 br_1_7 br_1_8 bl_0_10 br_1_10 bl_0_11
+ bl_1_11 br_0_11 br_1_11 bl_1_12 br_1_12 bl_0_13 bl_1_13 br_1_13 bl_1_14 br_0_14
+ br_1_14 bl_1_15 br_1_15 bl_1_16 br_1_16 br_1_17 bl_1_18 bl_1_19 br_0_19 br_1_19
+ bl_0_20 bl_1_20 br_0_20 br_1_20 br_1_21 br_0_22 br_1_22 bl_1_23 br_1_23 bl_1_24
+ br_1_24 bl_0_25 br_1_25 bl_1_27 br_1_27 bl_0_28 bl_1_28 br_1_28 bl_1_29 br_1_30
+ bl_0_31 br_1_31 vdd_uq0 vdd_uq1 vdd_uq2 vdd_uq3 vdd_uq4 vdd_uq5 vdd_uq6 vdd_uq7
+ vdd_uq8 vdd_uq10 vdd_uq13 vdd_uq22 sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_0/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_20/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_38_n79#
+ br_0_17 sky130_fd_bd_sram__openram_dp_cell_dummy_30/w_144_n79# bl_1_31 sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_400_n79# vdd_uq19 sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_400_n79#
+ br_0_25 sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_11/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_1/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_21/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_31/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_400_n79#
+ br_0_28 sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_38_n79#
+ bl_0_16 sky130_fd_bd_sram__openram_dp_cell_dummy_12/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_2/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_22/w_144_n79# vdd_uq17 vdd_uq26 bl_0_24
+ bl_1_1 sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_400_n79#
+ br_0_31 sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_400_n79#
+ bl_0_19 br_0_13 br_0_4 sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_13/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_3/w_144_n79# vdd_uq14 vdd_uq23 sky130_fd_bd_sram__openram_dp_cell_dummy_23/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_38_n79# bl_0_27 sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_38_n79#
+ br_0_8 br_0_16 sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_400_n79# br_0_7 bl_1_30
+ sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/w_144_n79#
+ vdd_uq20 vdd_uq11 sky130_fd_bd_sram__openram_dp_cell_dummy_4/w_144_n79# vdd_uq29
+ bl_1_3 sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_38_n79# bl_0_30 sky130_fd_bd_sram__openram_dp_cell_dummy_24/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_38_n79# br_0_24 bl_0_12 bl_0_3 sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_38_n79#
+ br_0_10 br_0_1 sky130_fd_bd_sram__openram_dp_cell_dummy_15/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/w_144_n79#
+ br_0_27 sky130_fd_bd_sram__openram_dp_cell_dummy_25/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_38_n79#
+ bl_0_15 sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_38_n79# bl_0_6 vdd sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_400_n79# vdd_uq18 sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_38_n79#
+ vdd_uq27 sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_400_n79# bl_0_23 bl_1_10
+ bl_1_0 sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_6/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_400_n79#
+ br_0_30 bl_0_18 bl_0_0 sky130_fd_bd_sram__openram_dp_cell_dummy_26/w_144_n79# br_0_12
+ br_0_3 sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_38_n79# vdd_uq15 vdd_uq24 sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_38_n79#
+ bl_0_26 bl_1_21 sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_7/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_400_n79#
+ bl_0_21 br_0_15 br_0_6 sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/w_144_n79#
+ vdd_uq12 vdd_uq30 vdd_uq21 bl_1_2 sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_400_n79# bl_0_29 br_0_23 br_1_18 br_1_9
+ sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_400_n79# bl_0_2 sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_18/w_144_n79# br_0_18 br_0_9 sky130_fd_bd_sram__openram_dp_cell_dummy_8/w_144_n79#
+ br_0_0 br_1_26 sky130_fd_bd_sram__openram_dp_cell_dummy_28/w_144_n79# vdd_uq9 sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_38_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_400_n79# br_0_26 sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_38_n79# bl_0_14 bl_0_5 sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_400_n79#
+ br_0_21 bl_1_22 sky130_fd_bd_sram__openram_dp_cell_dummy_19/w_144_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/w_144_n79#
+ vdd_uq28 br_1_29 bl_1_9 bl_0_22 sky130_fd_bd_sram__openram_dp_cell_dummy_29/w_144_n79#
+ bl_1_17 bl_1_8 sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_38_n79# br_1_2 br_0_29
+ bl_0_9 sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_400_n79#
+ bl_0_8 bl_0_17 sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_38_n79#
+ br_0_2 bl_1_26 wl_1_0 bl_1_25 sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_400_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_38_n79# vdd_uq16 vdd_uq25 gnd wl_0_0
Xsky130_fd_bd_sram__openram_dp_cell_dummy_30 gnd bl_0_1 br_0_1 bl_1_1 br_1_1 wl_0_0
+ wl_1_0 vdd_uq29 sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_30/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_30/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_10 gnd bl_0_21 br_0_21 bl_1_21 br_1_21 wl_0_0
+ wl_1_0 vdd_uq9 sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_10/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_10/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_20 gnd bl_0_11 br_0_11 bl_1_11 br_1_11 wl_0_0
+ wl_1_0 vdd_uq19 sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_20/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_20/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_21 gnd bl_0_10 br_0_10 bl_1_10 br_1_10 wl_0_0
+ wl_1_0 vdd_uq20 sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_21/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_21/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_31 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_0
+ wl_1_0 vdd_uq30 sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_31/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_31/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_11 gnd bl_0_20 br_0_20 bl_1_20 br_1_20 wl_0_0
+ wl_1_0 vdd_uq10 sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_11/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_11/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_22 gnd bl_0_9 br_0_9 bl_1_9 br_1_9 wl_0_0
+ wl_1_0 vdd_uq21 sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_22/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_22/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 gnd bl_0_31 br_0_31 bl_1_31 br_1_31 wl_0_0
+ wl_1_0 vdd_uq0 sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_0/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_0/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_12 gnd bl_0_19 br_0_19 bl_1_19 br_1_19 wl_0_0
+ wl_1_0 vdd_uq11 sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_12/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_12/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_23 gnd bl_0_8 br_0_8 bl_1_8 br_1_8 wl_0_0
+ wl_1_0 vdd_uq22 sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_23/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_23/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_1 gnd bl_0_30 br_0_30 bl_1_30 br_1_30 wl_0_0
+ wl_1_0 vdd sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_1/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_1/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_13 gnd bl_0_18 br_0_18 bl_1_18 br_1_18 wl_0_0
+ wl_1_0 vdd_uq12 sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_13/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_13/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_24 gnd bl_0_7 br_0_7 bl_1_7 br_1_7 wl_0_0
+ wl_1_0 vdd_uq23 sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_24/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_24/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_2 gnd bl_0_29 br_0_29 bl_1_29 br_1_29 wl_0_0
+ wl_1_0 vdd_uq1 sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_2/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_2/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_14 gnd bl_0_17 br_0_17 bl_1_17 br_1_17 wl_0_0
+ wl_1_0 vdd_uq13 sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_14/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_14/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_25 gnd bl_0_6 br_0_6 bl_1_6 br_1_6 wl_0_0
+ wl_1_0 vdd_uq24 sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_25/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_25/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_3 gnd bl_0_28 br_0_28 bl_1_28 br_1_28 wl_0_0
+ wl_1_0 vdd_uq2 sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_3/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_3/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_15 gnd bl_0_16 br_0_16 bl_1_16 br_1_16 wl_0_0
+ wl_1_0 vdd_uq14 sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_15/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_15/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_26 gnd bl_0_5 br_0_5 bl_1_5 br_1_5 wl_0_0
+ wl_1_0 vdd_uq25 sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_26/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_26/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_4 gnd bl_0_27 br_0_27 bl_1_27 br_1_27 wl_0_0
+ wl_1_0 vdd_uq3 sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_4/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_4/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_16 gnd bl_0_15 br_0_15 bl_1_15 br_1_15 wl_0_0
+ wl_1_0 vdd_uq15 sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_16/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_16/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_27 gnd bl_0_4 br_0_4 bl_1_4 br_1_4 wl_0_0
+ wl_1_0 vdd_uq26 sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_27/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_27/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_5 gnd bl_0_26 br_0_26 bl_1_26 br_1_26 wl_0_0
+ wl_1_0 vdd_uq4 sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_5/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_5/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_6 gnd bl_0_25 br_0_25 bl_1_25 br_1_25 wl_0_0
+ wl_1_0 vdd_uq5 sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_6/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_6/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_17 gnd bl_0_14 br_0_14 bl_1_14 br_1_14 wl_0_0
+ wl_1_0 vdd_uq16 sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_17/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_17/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_28 gnd bl_0_3 br_0_3 bl_1_3 br_1_3 wl_0_0
+ wl_1_0 vdd_uq27 sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_28/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_28/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_7 gnd bl_0_24 br_0_24 bl_1_24 br_1_24 wl_0_0
+ wl_1_0 vdd_uq6 sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_7/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_7/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_18 gnd bl_0_13 br_0_13 bl_1_13 br_1_13 wl_0_0
+ wl_1_0 vdd_uq17 sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_18/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_18/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_19 gnd bl_0_12 br_0_12 bl_1_12 br_1_12 wl_0_0
+ wl_1_0 vdd_uq18 sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_19/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_19/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_29 gnd bl_0_2 br_0_2 bl_1_2 br_1_2 wl_0_0
+ wl_1_0 vdd_uq28 sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_29/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_29/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_8 gnd bl_0_23 br_0_23 bl_1_23 br_1_23 wl_0_0
+ wl_1_0 vdd_uq7 sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_8/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_8/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_dummy_9 gnd bl_0_22 br_0_22 bl_1_22 br_1_22 wl_0_0
+ wl_1_0 vdd_uq8 sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_38_n79# sky130_fd_bd_sram__openram_dp_cell_dummy_9/w_144_n79#
+ sky130_fd_bd_sram__openram_dp_cell_dummy_9/a_400_n79# sky130_fd_bd_sram__openram_dp_cell_dummy
.ends

.subckt sky130_fd_bd_sram__openram_dp_cell_replica gnd bl0 br0 bl1 br1 wl0 wl1 vdd
+ a_38_n79# a_400_n79#
X0 gnd gnd bl1 gnd sky130_fd_pr__special_nfet_latch ad=1.0032p pd=13.14u as=0.0504p ps=0.9u w=0.21u l=0.08u
X1 a_38_133# wl0 a_38_133# vdd sky130_fd_pr__special_pfet_pass ad=0.035p pd=0.78u as=0p ps=0u w=0.07u l=0.15u
X2 vdd wl1 br1 gnd sky130_fd_pr__special_nfet_latch ad=0.3088p pd=4.43u as=0.0504p ps=0.9u w=0.21u l=0.15u
X3 gnd gnd a_400_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X4 vdd a_38_133# gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.2768p ps=4u w=0.21u l=0.15u
X5 vdd wl1 vdd vdd sky130_fd_pr__special_pfet_pass ad=0.0714p pd=1.58u as=0p ps=0u w=0.07u l=0.15u
X6 a_38_133# wl1 bl1 gnd sky130_fd_pr__special_nfet_latch ad=0.3463p pd=4.93u as=0p ps=0u w=0.21u l=0.15u
X7 gnd gnd a_38_n79# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.0252p ps=0.66u w=0.21u l=0.08u
X8 gnd gnd br1 gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.08u
X9 a_38_133# vdd gnd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X10 br0 wl0 vdd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.1974p ps=3.44u w=0.21u l=0.15u
X11 gnd a_38_133# vdd gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
X12 a_38_133# vdd vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=0.14u l=0.15u
X13 vdd a_38_133# vdd vdd sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=0.14u l=0.15u
X14 bl0 wl0 a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0.105p ps=1.84u w=0.21u l=0.15u
X15 gnd vdd a_38_133# gnd sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=0.21u l=0.15u
.ends

.subckt subbyte2_replica_column wl_0_1 wl_1_1 wl_0_2 wl_1_2 wl_0_3 wl_0_4 wl_0_5 wl_1_5
+ wl_0_6 wl_0_7 wl_0_8 wl_1_8 wl_1_10 wl_1_11 wl_1_13 wl_1_14 wl_0_15 wl_0_16 wl_1_16
+ wl_0_17 wl_1_17 wl_0_18 wl_0_19 wl_1_19 wl_1_20 wl_1_22 wl_1_23 wl_1_25 wl_0_26
+ wl_1_26 wl_0_27 wl_0_28 wl_1_28 wl_0_29 wl_1_29 wl_1_32 wl_1_34 wl_1_35 wl_0_37
+ wl_0_38 wl_1_38 wl_0_39 wl_1_40 wl_1_41 wl_1_43 wl_1_44 wl_1_46 wl_1_47 wl_0_48
+ wl_0_49 wl_1_49 wl_1_50 wl_1_52 wl_1_53 wl_0_54 wl_1_54 wl_1_55 wl_1_57 wl_1_58
+ wl_0_59 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63 wl_1_64 wl_1_65 wl_0_35 wl_0_47
+ wl_0_20 wl_0_11 wl_0_55 wl_0_41 wl_0_32 wl_0_23 wl_0_14 wl_0_58 wl_0_53 wl_0_44
+ wl_1_7 wl_0_62 wl_0_61 wl_0_25 wl_0_46 wl_0_64 wl_0_10 wl_1_4 wl_0_50 wl_0_40 wl_0_31
+ wl_0_13 wl_0_65 wl_0_22 wl_0_57 wl_0_52 wl_0_43 wl_0_34 wl_1_15 wl_1_6 wl_0_60 wl_1_37
+ wl_1_45 wl_1_36 wl_1_27 wl_1_18 wl_1_0 wl_1_9 wl_0_63 wl_0_45 wl_0_36 wl_0_9 wl_0_0
+ wl_1_31 wl_1_48 wl_1_39 wl_1_21 wl_1_30 wl_1_12 wl_1_3 wl_0_30 wl_0_21 wl_0_12 wl_1_56
+ wl_1_51 wl_1_42 br_0_0 wl_1_33 wl_1_24 wl_0_56 vdd wl_0_51 wl_0_42 wl_0_33 wl_0_24
+ bl_1_0 br_1_0 bl_0_0 gnd
Xsky130_fd_bd_sram__openram_dp_cell_replica_50 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_14
+ wl_1_14 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_60 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_4
+ wl_1_4 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_61 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_3
+ wl_1_3 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_40 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_24
+ wl_1_24 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_51 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_13
+ wl_1_13 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_62 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_2
+ wl_1_2 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_30 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_34
+ wl_1_34 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_41 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_23
+ wl_1_23 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_52 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_12
+ wl_1_12 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_63 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_1
+ wl_1_1 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_65
+ wl_1_65 vdd bl_1_0 vdd br_1_0 sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_replica_20 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_44
+ wl_1_44 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_31 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_33
+ wl_1_33 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_42 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_22
+ wl_1_22 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_53 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_11
+ wl_1_11 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_64 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_0
+ wl_1_0 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_10 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_54
+ wl_1_54 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_21 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_43
+ wl_1_43 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_32 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_32
+ wl_1_32 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_43 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_21
+ wl_1_21 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_54 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_10
+ wl_1_10 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_11 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_53
+ wl_1_53 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_22 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_42
+ wl_1_42 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_33 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_31
+ wl_1_31 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_44 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_20
+ wl_1_20 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_55 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_9
+ wl_1_9 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_12 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_52
+ wl_1_52 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_23 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_41
+ wl_1_41 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_34 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_30
+ wl_1_30 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_45 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_19
+ wl_1_19 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_56 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_8
+ wl_1_8 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_13 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_51
+ wl_1_51 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_24 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_40
+ wl_1_40 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_35 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_29
+ wl_1_29 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_46 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_18
+ wl_1_18 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_57 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_7
+ wl_1_7 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_0 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_64
+ wl_1_64 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_14 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_50
+ wl_1_50 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_15 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_49
+ wl_1_49 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_25 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_39
+ wl_1_39 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_26 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_38
+ wl_1_38 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_36 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_28
+ wl_1_28 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_37 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_27
+ wl_1_27 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_47 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_17
+ wl_1_17 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_48 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_16
+ wl_1_16 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_58 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_6
+ wl_1_6 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_59 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_5
+ wl_1_5 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_1 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_63
+ wl_1_63 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_16 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_48
+ wl_1_48 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_27 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_37
+ wl_1_37 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_38 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_26
+ wl_1_26 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_49 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_15
+ wl_1_15 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_2 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_62
+ wl_1_62 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_17 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_47
+ wl_1_47 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_28 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_36
+ wl_1_36 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_39 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_25
+ wl_1_25 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_3 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_61
+ wl_1_61 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_18 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_46
+ wl_1_46 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_29 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_35
+ wl_1_35 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_4 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_60
+ wl_1_60 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_19 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_45
+ wl_1_45 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_5 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_59
+ wl_1_59 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_6 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_58
+ wl_1_58 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_7 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_57
+ wl_1_57 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_8 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_56
+ wl_1_56 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_9 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_55
+ wl_1_55 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
.ends

.subckt subbyte2_replica_column_0 wl_1_0 wl_0_1 wl_0_2 wl_1_2 wl_0_3 wl_1_3 wl_0_4
+ wl_0_5 wl_0_6 wl_1_6 wl_0_7 wl_0_8 wl_0_9 wl_1_9 wl_1_10 wl_1_11 wl_1_12 wl_1_14
+ wl_0_15 wl_1_15 wl_0_16 wl_0_17 wl_1_17 wl_0_18 wl_1_18 wl_0_19 wl_1_20 wl_1_21
+ wl_1_23 wl_1_24 wl_0_26 wl_0_27 wl_1_27 wl_0_28 wl_0_29 wl_1_29 wl_1_30 wl_1_32
+ wl_1_33 wl_1_35 wl_1_36 wl_0_37 wl_0_38 wl_1_38 wl_0_39 wl_1_39 wl_1_40 wl_1_41
+ wl_1_42 wl_1_44 wl_1_45 wl_1_47 wl_0_48 wl_1_48 wl_0_49 wl_1_50 wl_1_51 wl_1_53
+ wl_1_54 wl_0_55 wl_1_55 wl_1_56 wl_1_58 wl_0_59 wl_1_59 wl_0_60 wl_1_60 wl_1_61
+ wl_1_62 wl_0_63 wl_1_63 wl_1_64 wl_1_65 wl_0_36 wl_0_30 wl_0_21 wl_0_12 wl_0_51
+ wl_0_42 wl_0_33 wl_0_24 wl_0_54 wl_0_45 wl_1_8 wl_0_65 wl_0_47 wl_0_20 wl_0_11 wl_1_5
+ wl_0_56 wl_0_41 wl_0_32 wl_0_14 wl_0_0 wl_0_23 wl_0_58 wl_0_44 wl_0_53 wl_0_35 wl_1_26
+ wl_1_16 wl_1_7 wl_0_62 wl_0_61 wl_1_46 wl_1_37 wl_1_28 wl_1_19 wl_1_1 wl_0_46 wl_0_64
+ wl_0_10 wl_1_49 wl_1_22 wl_1_31 wl_1_13 wl_1_4 wl_0_50 wl_0_40 wl_0_31 wl_0_13 wl_0_22
+ wl_1_57 wl_1_52 wl_1_43 br_0_0 wl_1_34 wl_1_25 wl_0_57 vdd wl_0_52 wl_0_43 wl_0_34
+ wl_0_25 bl_1_0 br_1_0 bl_0_0 gnd
Xsky130_fd_bd_sram__openram_dp_cell_replica_50 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_15
+ wl_1_15 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_60 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_5
+ wl_1_5 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_61 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_4
+ wl_1_4 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_40 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_25
+ wl_1_25 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_51 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_14
+ wl_1_14 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_62 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_3
+ wl_1_3 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_30 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_35
+ wl_1_35 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_41 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_24
+ wl_1_24 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_52 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_13
+ wl_1_13 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_63 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_2
+ wl_1_2 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_20 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_45
+ wl_1_45 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_31 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_34
+ wl_1_34 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_42 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_23
+ wl_1_23 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_53 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_12
+ wl_1_12 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_64 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_1
+ wl_1_1 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_dummy_0 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_0
+ wl_1_0 vdd bl_1_0 vdd br_1_0 sky130_fd_bd_sram__openram_dp_cell_dummy
Xsky130_fd_bd_sram__openram_dp_cell_replica_10 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_55
+ wl_1_55 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_21 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_44
+ wl_1_44 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_32 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_33
+ wl_1_33 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_43 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_22
+ wl_1_22 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_54 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_11
+ wl_1_11 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_11 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_54
+ wl_1_54 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_22 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_43
+ wl_1_43 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_33 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_32
+ wl_1_32 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_44 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_21
+ wl_1_21 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_55 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_10
+ wl_1_10 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_12 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_53
+ wl_1_53 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_23 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_42
+ wl_1_42 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_34 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_31
+ wl_1_31 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_45 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_20
+ wl_1_20 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_56 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_9
+ wl_1_9 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_13 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_52
+ wl_1_52 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_24 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_41
+ wl_1_41 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_35 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_30
+ wl_1_30 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_46 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_19
+ wl_1_19 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_57 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_8
+ wl_1_8 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_0 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_65
+ wl_1_65 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_14 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_51
+ wl_1_51 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_15 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_50
+ wl_1_50 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_25 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_40
+ wl_1_40 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_26 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_39
+ wl_1_39 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_36 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_29
+ wl_1_29 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_37 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_28
+ wl_1_28 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_47 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_18
+ wl_1_18 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_48 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_17
+ wl_1_17 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_58 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_7
+ wl_1_7 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_59 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_6
+ wl_1_6 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_1 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_64
+ wl_1_64 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_16 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_49
+ wl_1_49 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_27 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_38
+ wl_1_38 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_38 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_27
+ wl_1_27 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_49 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_16
+ wl_1_16 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_2 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_63
+ wl_1_63 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_17 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_48
+ wl_1_48 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_28 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_37
+ wl_1_37 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_39 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_26
+ wl_1_26 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_3 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_62
+ wl_1_62 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_18 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_47
+ wl_1_47 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_29 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_36
+ wl_1_36 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_4 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_61
+ wl_1_61 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_19 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_46
+ wl_1_46 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_5 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_60
+ wl_1_60 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_6 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_59
+ wl_1_59 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_7 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_58
+ wl_1_58 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_8 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_57
+ wl_1_57 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
Xsky130_fd_bd_sram__openram_dp_cell_replica_9 gnd bl_0_0 br_0_0 bl_1_0 br_1_0 wl_0_56
+ wl_1_56 vdd bl_1_0 br_1_0 sky130_fd_bd_sram__openram_dp_cell_replica
.ends

.subckt subbyte2_replica_bitcell_array bl_1_12 br_0_19 bl_1_23 wl_0_1 wl_0_2 wl_0_15
+ wl_0_16 wl_0_17 wl_0_26 wl_0_28 wl_0_37 wl_0_48 wl_0_59 vdd_uq98 vdd_uq6 vdd_uq7
+ vdd_uq85 vdd_uq96 vdd_uq97 vdd_uq5 vdd_uq84 vdd_uq95 vdd_uq4 vdd_uq83 vdd_uq94 vdd_uq3
+ vdd_uq9 vdd_uq78 vdd_uq86 vdd_uq87 vdd_uq88 vdd_uq2 vdd_uq89 wl_1_44 wl_1_35 wl_1_26
+ br_1_24 bl_0_11 br_1_28 br_0_1 bl_0_22 wl_0_8 bl_0_7 bl_0_18 wl_0_35 bl_1_17 wl_0_63
+ wl_0_46 bl_1_6 wl_0_7 rbl_br_1_0 wl_0_19 bl_0_10 bl_0_21 br_0_4 wl_0_60 br_1_3 bl_1_9
+ br_0_25 wl_1_56 vdd_uq66 rbl_bl_1_1 wl_1_33 wl_1_30 br_1_31 wl_1_24 wl_1_21 br_0_14
+ vdd_uq91 rbl_wl_1_1 vdd vdd_uq90 wl_1_15 bl_1_16 vdd_uq79 wl_1_12 br_1_6 rbl_br_1_1
+ vdd_uq99 br_1_20 bl_1_26 bl_1_15 wl_0_57 br_0_24 wl_0_62 wl_0_51 br_1_16 br_1_27
+ br_1_13 bl_0_3 br_1_12 wl_0_45 br_1_23 bl_1_29 bl_0_17 wl_0_13 bl_0_6 br_0_29 br_0_18
+ wl_0_54 bl_1_2 vdd_uq1 vdd_uq93 vdd_uq82 wl_1_53 rbl_br_0_0 bl_1_0 bl_0_5 bl_1_1
+ rbl_wl_0_1 wl_1_50 wl_0_27 br_1_15 wl_0_10 wl_1_41 br_0_3 bl_0_9 br_1_26 wl_0_18
+ bl_1_5 bl_0_20 wl_1_47 br_0_0 br_1_2 bl_1_8 bl_0_31 bl_1_19 wl_0_9 bl_1_20 bl_1_4
+ bl_1_31 wl_0_56 wl_0_0 wl_0_42 bl_1_3 rbl_bl_0_1 br_1_29 bl_0_8 rbl_bl_0_0 wl_0_30
+ wl_0_38 br_0_31 wl_1_45 br_0_2 wl_0_24 wl_1_38 br_0_10 wl_0_21 wl_0_29 br_0_21 bl_0_27
+ wl_1_36 bl_0_23 rbl_wl_1_0 wl_1_32 wl_1_29 bl_0_16 wl_0_12 br_0_6 bl_0_12 rbl_br_0_1
+ wl_1_27 wl_1_23 bl_0_14 wl_0_6 wl_1_20 bl_0_25 bl_1_22 wl_0_3 br_1_5 br_0_20 bl_0_26
+ wl_1_18 wl_1_6 br_1_9 br_0_8 vdd_uq8 wl_1_3 bl_1_11 wl_1_11 br_1_1 bl_1_7 br_0_9
+ bl_0_15 bl_1_18 wl_1_28 wl_1_9 bl_1_30 wl_1_61 wl_0_61 wl_1_58 wl_0_39 wl_0_52 wl_1_2
+ wl_0_41 br_1_0 br_0_5 wl_0_49 bl_0_30 br_0_16 wl_1_19 wl_1_0 wl_1_52 br_0_27 wl_1_49
+ wl_0_43 wl_1_57 br_0_13 wl_0_32 wl_0_40 wl_1_10 wl_1_43 br_0_12 wl_0_20 wl_0_55
+ wl_0_44 wl_0_33 wl_0_22 vdd_uq0 wl_0_11 vdd_uq80 wl_1_40 br_0_23 bl_0_29 br_1_4
+ wl_0_34 wl_0_23 wl_0_31 bl_1_13 br_1_22 wl_1_1 wl_1_46 wl_1_34 br_1_18 bl_1_24 wl_1_42
+ wl_1_31 bl_0_28 wl_1_39 br_1_19 bl_1_25 wl_1_55 wl_0_4 br_1_7 wl_1_17 wl_1_37 br_0_28
+ wl_1_25 br_0_11 br_0_17 br_1_17 wl_1_14 wl_0_58 wl_0_47 br_1_8 wl_0_36 bl_1_14 wl_0_25
+ wl_0_14 wl_1_22 br_0_22 wl_0_5 bl_0_2 wl_1_8 wl_1_16 wl_1_5 wl_1_13 bl_1_28 vdd_uq92
+ vdd_uq81 wl_1_63 bl_1_21 bl_1_10 wl_1_7 wl_0_53 bl_0_0 br_1_11 wl_1_60 bl_0_24 bl_0_13
+ wl_1_4 br_0_7 bl_0_1 br_1_10 wl_1_48 br_1_25 wl_1_54 br_0_15 br_1_21 bl_0_4 bl_1_27
+ br_0_30 bl_0_19 wl_1_62 wl_0_50 br_1_30 rbl_wl_0_0 br_0_26 wl_1_51 wl_1_59 rbl_bl_1_0
+ br_1_14 gnd
Xsubbyte2_bitcell_array_0 bl_1_12 br_0_19 bl_1_23 wl_0_2 wl_0_15 wl_0_16 wl_0_17 wl_0_26
+ wl_0_37 wl_0_38 wl_0_48 wl_0_49 wl_1_53 wl_1_62 wl_1_63 vdd_uq6 vdd_uq9 vdd_uq81
+ vdd_uq82 vdd_uq83 vdd_uq87 vdd_uq88 vdd_uq93 vdd_uq98 bl_1_25 bl_1_10 br_1_31 br_1_16
+ br_1_15 bl_1_22 bl_1_18 bl_1_7 bl_1_3 br_1_20 br_1_9 bl_1_0 bl_1_12 bl_1_26 bl_1_0
+ bl_1_16 br_1_8 br_1_26 br_1_19 br_1_8 bl_1_28 bl_1_13 bl_1_27 bl_1_9 br_1_30 br_1_12
+ br_1_7 bl_1_30 bl_1_24 bl_1_20 bl_1_9 br_1_19 br_1_1 bl_1_5 bl_1_24 br_1_29 bl_1_17
+ bl_1_2 br_1_23 bl_1_7 bl_1_21 br_1_18 br_1_0 bl_1_6 bl_1_31 bl_1_26 bl_1_15 bl_1_11
+ br_1_22 br_1_11 br_1_22 br_1_11 br_1_6 bl_1_8 bl_1_22 bl_1_4 br_1_15 br_1_10 br_1_10
+ bl_1_19 bl_1_4 br_1_4 bl_1_23 bl_1_19 br_1_14 br_1_31 br_1_9 bl_1_28 br_1_26 bl_1_13
+ br_1_21 br_1_3 bl_1_16 br_1_21 br_1_3 bl_1_1 bl_1_25 bl_1_10 bl_1_6 br_1_25 br_1_14
+ br_1_7 br_1_30 br_1_2 bl_1_15 br_1_25 br_1_20 br_1_2 bl_1_3 bl_1_17 bl_1_2 br_1_13
+ br_1_24 br_1_13 bl_1_21 br_1_0 bl_1_30 br_1_18 bl_1_18 wl_0_25 br_1_12 bl_1_27 bl_1_23
+ bl_1_12 br_1_29 bl_1_8 br_1_24 wl_1_8 br_1_17 br_1_6 wl_0_53 br_1_17 wl_0_8 br_1_1
+ wl_1_16 wl_0_63 wl_1_7 bl_1_5 bl_1_1 wl_0_7 wl_0_62 br_1_28 bl_1_14 br_1_5 wl_1_44
+ wl_1_35 br_1_28 br_1_23 br_1_5 wl_0_44 wl_0_29 bl_0_21 bl_1_29 bl_0_1 wl_0_35 br_1_31
+ wl_1_28 br_0_18 bl_0_4 wl_1_11 vdd_uq2 vdd_uq90 wl_0_58 bl_1_20 wl_1_2 wl_1_57 br_0_25
+ br_0_5 bl_0_11 br_0_1 bl_0_7 br_1_17 wl_1_22 bl_1_14 wl_1_13 bl_1_26 br_1_20 bl_1_6
+ br_0_24 vdd_uq84 bl_0_10 wl_0_5 br_0_4 wl_0_60 wl_1_54 br_1_23 bl_1_29 br_1_3 bl_1_9
+ bl_0_17 vdd_uq97 bl_0_31 br_0_7 bl_0_30 wl_1_42 wl_0_46 wl_1_19 wl_1_33 vdd_uq5
+ br_1_27 br_1_16 wl_1_45 br_0_31 wl_1_24 br_1_30 br_1_10 vdd_uq94 wl_0_20 vdd_uq78
+ wl_0_28 bl_0_24 br_0_14 wl_1_36 wl_0_11 bl_1_16 br_1_26 wl_0_19 br_1_6 bl_0_0 bl_0_20
+ wl_1_27 bl_1_19 wl_1_18 wl_1_10 br_1_29 br_1_9 bl_1_15 wl_0_57 wl_1_9 wl_1_1 wl_0_40
+ vdd_uq95 br_1_16 wl_1_0 wl_1_48 br_1_13 wl_1_56 wl_0_31 bl_0_2 br_0_17 bl_0_23 bl_0_3
+ br_1_12 wl_1_55 wl_1_39 vdd_uq91 vdd_uq3 wl_0_22 br_0_21 bl_0_27 wl_1_46 wl_1_30
+ wl_1_38 wl_1_25 wl_0_13 bl_0_26 br_0_20 bl_0_6 br_1_11 wl_1_37 wl_1_21 bl_0_25 wl_1_29
+ bl_1_2 bl_1_22 bl_1_18 wl_1_4 wl_1_12 wl_0_51 bl_1_20 bl_1_0 wl_1_59 wl_1_3 bl_0_5
+ bl_1_1 bl_1_21 vdd_uq85 vdd_uq89 wl_0_30 br_0_27 bl_0_13 wl_1_50 br_1_27 br_1_15
+ wl_0_21 wl_0_54 br_0_23 br_0_3 wl_1_41 bl_0_29 bl_0_9 br_1_19 bl_1_25 bl_1_5 vdd
+ wl_1_47 br_0_0 br_1_22 bl_1_28 br_1_2 bl_1_8 wl_0_4 br_1_14 bl_1_24 wl_0_12 bl_0_28
+ wl_1_20 br_1_18 bl_1_4 wl_1_15 wl_0_3 br_0_22 wl_0_42 wl_0_50 bl_1_3 bl_0_8 wl_1_58
+ wl_0_33 vdd_uq86 wl_0_41 br_0_2 wl_0_45 vdd_uq1 wl_1_49 wl_0_24 wl_0_32 br_0_30
+ br_0_10 wl_0_36 wl_1_32 br_0_28 vdd_uq7 wl_1_40 bl_1_27 br_1_4 wl_0_23 bl_0_16 br_0_6
+ bl_0_12 br_0_26 wl_0_27 wl_1_23 bl_0_14 vdd_uq79 wl_1_31 br_1_5 br_1_25 wl_0_6 br_1_21
+ wl_1_26 wl_0_14 bl_0_19 wl_1_6 wl_0_18 br_0_8 wl_1_14 bl_1_11 wl_0_10 wl_0_61 wl_1_17
+ br_1_1 bl_1_7 br_0_29 br_0_9 bl_0_15 wl_1_61 wl_0_9 wl_1_5 wl_0_1 wl_0_52 br_1_0
+ bl_1_29 br_0_16 wl_1_52 wl_0_0 wl_1_60 bl_1_11 vdd_uq80 wl_0_56 wl_0_43 br_0_13
+ br_1_27 vdd_uq99 wl_0_59 bl_1_31 br_0_12 wl_1_43 vdd_uq8 wl_0_55 br_1_28 bl_1_17
+ wl_0_39 wl_1_51 bl_1_14 br_1_8 vdd_uq96 br_1_24 br_1_4 wl_0_47 bl_1_10 wl_0_34 bl_1_30
+ bl_0_22 bl_0_18 br_1_7 bl_1_13 gnd br_0_15 vdd_uq92 br_0_11 wl_1_34 bl_1_31 vdd_uq4
+ subbyte2_bitcell_array
Xsubbyte2_dummy_array_0 br_1_0 bl_0_1 br_1_1 br_1_3 bl_0_4 bl_1_4 br_1_4 bl_1_5 br_0_5
+ br_1_5 bl_1_6 br_1_6 bl_0_7 bl_1_7 br_1_7 br_1_8 bl_0_10 br_1_10 bl_0_11 bl_1_11
+ br_0_11 br_1_11 bl_1_12 br_1_12 bl_0_13 bl_1_13 br_1_13 bl_1_14 br_0_14 br_1_14
+ bl_1_15 br_1_15 bl_1_16 br_1_16 br_1_17 bl_1_18 bl_1_19 br_0_19 br_1_19 bl_0_20
+ bl_1_20 br_0_20 br_1_20 br_1_21 br_0_22 br_1_22 bl_1_23 br_1_23 bl_1_24 br_1_24
+ bl_0_25 br_1_25 bl_1_27 br_1_27 bl_0_28 bl_1_28 br_1_28 bl_1_29 br_1_30 bl_0_31
+ br_1_31 vdd vdd_uq2 vdd_uq3 vdd_uq4 vdd_uq5 vdd_uq6 vdd_uq7 vdd_uq8 vdd_uq9 vdd_uq79
+ vdd_uq82 vdd_uq91 bl_1_31 br_1_16 br_1_26 br_1_6 bl_1_14 vdd_uq78 vdd vdd_uq88 bl_1_18
+ br_0_17 vdd_uq98 bl_1_31 br_1_15 br_1_25 vdd_uq88 br_1_5 br_0_25 bl_1_4 vdd_uq79
+ vdd_uq1 bl_1_22 vdd_uq89 bl_1_8 vdd_uq99 bl_1_26 br_1_14 br_1_24 br_0_28 br_1_4
+ bl_1_30 bl_0_16 vdd_uq80 vdd_uq2 vdd_uq90 vdd_uq86 vdd_uq95 bl_0_24 bl_1_1 br_1_13
+ br_1_23 br_0_31 bl_1_13 br_1_3 bl_0_19 br_0_13 br_0_4 bl_1_17 vdd_uq81 vdd_uq3 vdd_uq83
+ vdd_uq92 vdd_uq91 bl_1_21 bl_0_27 br_1_12 br_1_22 bl_1_3 br_0_8 br_0_16 br_1_2 br_0_7
+ bl_1_30 bl_1_7 vdd_uq82 vdd_uq89 vdd_uq80 vdd_uq4 vdd_uq98 bl_1_3 bl_1_25 bl_0_30
+ vdd_uq92 bl_1_11 br_0_24 bl_0_12 bl_0_3 bl_1_29 br_0_10 br_0_1 vdd_uq83 vdd_uq5
+ br_0_27 vdd_uq93 bl_1_1 bl_0_15 bl_1_12 bl_0_6 vdd_uq1 br_1_21 br_1_31 vdd_uq87
+ bl_1_16 vdd_uq96 br_1_11 bl_0_23 bl_1_10 bl_1_0 bl_1_20 vdd_uq84 vdd_uq6 br_1_1
+ br_0_30 bl_0_18 bl_0_0 vdd_uq94 br_0_12 br_0_3 bl_1_2 vdd_uq84 vdd_uq93 br_1_20
+ br_1_30 bl_1_6 bl_0_26 bl_1_21 br_1_10 bl_1_24 bl_1_10 vdd_uq85 vdd_uq7 br_1_0 bl_0_21
+ br_0_15 br_0_6 bl_1_28 vdd_uq95 vdd_uq81 vdd_uq99 vdd_uq90 bl_1_2 br_1_19 br_1_29
+ bl_0_29 br_0_23 br_1_18 br_1_9 br_1_9 bl_0_2 bl_1_0 vdd_uq86 br_0_18 br_0_9 vdd_uq8
+ br_0_0 br_1_26 vdd_uq96 vdd_uq78 bl_1_15 br_1_18 br_0_26 br_1_28 bl_1_19 bl_0_14
+ bl_0_5 br_1_8 br_0_21 bl_1_22 vdd_uq87 vdd_uq9 vdd_uq97 br_1_29 bl_1_9 bl_0_22 vdd_uq97
+ bl_1_17 bl_1_8 bl_1_5 br_1_2 br_0_29 bl_0_9 bl_1_23 br_1_17 bl_0_8 bl_0_17 br_1_27
+ bl_1_9 br_0_2 bl_1_26 rbl_wl_1_1 bl_1_25 br_1_7 bl_1_27 vdd_uq85 vdd_uq94 gnd rbl_wl_1_0
+ subbyte2_dummy_array
Xsubbyte2_replica_column_0 wl_0_0 wl_1_0 wl_0_1 wl_1_1 wl_0_2 wl_0_3 wl_0_4 wl_1_4
+ wl_0_5 wl_0_6 wl_0_7 wl_1_7 wl_1_9 wl_1_10 wl_1_12 wl_1_13 wl_0_14 wl_0_15 wl_1_15
+ wl_0_16 wl_1_16 wl_0_17 wl_0_18 wl_1_18 wl_1_19 wl_1_21 wl_1_22 wl_1_24 wl_0_25
+ wl_1_25 wl_0_26 wl_0_27 wl_1_27 wl_0_28 wl_1_28 wl_1_31 wl_1_33 wl_1_34 wl_0_36
+ wl_0_37 wl_1_37 wl_0_38 wl_1_39 wl_1_40 wl_1_42 wl_1_43 wl_1_45 wl_1_46 wl_0_47
+ wl_0_48 wl_1_48 wl_1_49 wl_1_51 wl_1_52 wl_0_53 wl_1_53 wl_1_54 wl_1_56 wl_1_57
+ wl_0_58 wl_1_58 wl_1_59 wl_1_60 wl_1_61 wl_1_62 wl_1_63 rbl_wl_1_1 wl_0_34 wl_0_46
+ wl_0_19 wl_0_10 wl_0_54 wl_0_40 wl_0_31 wl_0_22 wl_0_13 wl_0_57 wl_0_52 wl_0_43
+ wl_1_6 wl_0_61 wl_0_60 wl_0_24 wl_0_45 wl_0_63 wl_0_9 wl_1_3 wl_0_49 wl_0_39 wl_0_30
+ wl_0_12 rbl_wl_1_0 wl_0_21 wl_0_56 wl_0_51 wl_0_42 wl_0_33 wl_1_14 wl_1_5 wl_0_59
+ wl_1_36 wl_1_44 wl_1_35 wl_1_26 wl_1_17 rbl_wl_0_1 wl_1_8 wl_0_62 wl_0_44 wl_0_35
+ wl_0_8 rbl_wl_0_0 wl_1_30 wl_1_47 wl_1_38 wl_1_20 wl_1_29 wl_1_11 wl_1_2 wl_0_29
+ wl_0_20 wl_0_11 wl_1_55 wl_1_50 wl_1_41 rbl_br_0_0 wl_1_32 wl_1_23 wl_0_55 vdd_uq66
+ wl_0_50 wl_0_41 wl_0_32 wl_0_23 rbl_bl_1_0 rbl_br_1_0 rbl_bl_0_0 gnd subbyte2_replica_column
Xsubbyte2_dummy_array_1 br_1_0 bl_0_1 br_1_1 br_1_3 bl_0_4 bl_1_4 br_1_4 bl_1_5 br_0_5
+ br_1_5 bl_1_6 br_1_6 bl_0_7 bl_1_7 br_1_7 br_1_8 bl_0_10 br_1_10 bl_0_11 bl_1_11
+ br_0_11 br_1_11 bl_1_12 br_1_12 bl_0_13 bl_1_13 br_1_13 bl_1_14 br_0_14 br_1_14
+ bl_1_15 br_1_15 bl_1_16 br_1_16 br_1_17 bl_1_18 bl_1_19 br_0_19 br_1_19 bl_0_20
+ bl_1_20 br_0_20 br_1_20 br_1_21 br_0_22 br_1_22 bl_1_23 br_1_23 bl_1_24 br_1_24
+ bl_0_25 br_1_25 bl_1_27 br_1_27 bl_0_28 bl_1_28 br_1_28 bl_1_29 br_1_30 bl_0_31
+ br_1_31 vdd vdd_uq2 vdd_uq3 vdd_uq4 vdd_uq5 vdd_uq6 vdd_uq7 vdd_uq8 vdd_uq9 vdd_uq79
+ vdd_uq82 vdd_uq91 bl_1_31 br_1_16 br_1_26 br_1_6 bl_1_14 vdd_uq78 vdd vdd_uq88 bl_1_18
+ br_0_17 vdd_uq98 bl_1_31 br_1_15 br_1_25 vdd_uq88 br_1_5 br_0_25 bl_1_4 vdd_uq79
+ vdd_uq1 bl_1_22 vdd_uq89 bl_1_8 vdd_uq99 bl_1_26 br_1_14 br_1_24 br_0_28 br_1_4
+ bl_1_30 bl_0_16 vdd_uq80 vdd_uq2 vdd_uq90 vdd_uq86 vdd_uq95 bl_0_24 bl_1_1 br_1_13
+ br_1_23 br_0_31 bl_1_13 br_1_3 bl_0_19 br_0_13 br_0_4 bl_1_17 vdd_uq81 vdd_uq3 vdd_uq83
+ vdd_uq92 vdd_uq91 bl_1_21 bl_0_27 br_1_12 br_1_22 bl_1_3 br_0_8 br_0_16 br_1_2 br_0_7
+ bl_1_30 bl_1_7 vdd_uq82 vdd_uq89 vdd_uq80 vdd_uq4 vdd_uq98 bl_1_3 bl_1_25 bl_0_30
+ vdd_uq92 bl_1_11 br_0_24 bl_0_12 bl_0_3 bl_1_29 br_0_10 br_0_1 vdd_uq83 vdd_uq5
+ br_0_27 vdd_uq93 bl_1_1 bl_0_15 bl_1_12 bl_0_6 vdd_uq1 br_1_21 br_1_31 vdd_uq87
+ bl_1_16 vdd_uq96 br_1_11 bl_0_23 bl_1_10 bl_1_0 bl_1_20 vdd_uq84 vdd_uq6 br_1_1
+ br_0_30 bl_0_18 bl_0_0 vdd_uq94 br_0_12 br_0_3 bl_1_2 vdd_uq84 vdd_uq93 br_1_20
+ br_1_30 bl_1_6 bl_0_26 bl_1_21 br_1_10 bl_1_24 bl_1_10 vdd_uq85 vdd_uq7 br_1_0 bl_0_21
+ br_0_15 br_0_6 bl_1_28 vdd_uq95 vdd_uq81 vdd_uq99 vdd_uq90 bl_1_2 br_1_19 br_1_29
+ bl_0_29 br_0_23 br_1_18 br_1_9 br_1_9 bl_0_2 bl_1_0 vdd_uq86 br_0_18 br_0_9 vdd_uq8
+ br_0_0 br_1_26 vdd_uq96 vdd_uq78 bl_1_15 br_1_18 br_0_26 br_1_28 bl_1_19 bl_0_14
+ bl_0_5 br_1_8 br_0_21 bl_1_22 vdd_uq87 vdd_uq9 vdd_uq97 br_1_29 bl_1_9 bl_0_22 vdd_uq97
+ bl_1_17 bl_1_8 bl_1_5 br_1_2 br_0_29 bl_0_9 bl_1_23 br_1_17 bl_0_8 bl_0_17 br_1_27
+ bl_1_9 br_0_2 bl_1_26 rbl_wl_0_1 bl_1_25 br_1_7 bl_1_27 vdd_uq85 vdd_uq94 gnd rbl_wl_0_0
+ subbyte2_dummy_array
Xsubbyte2_replica_column_0_0 rbl_wl_0_1 wl_0_0 wl_0_1 wl_1_1 wl_0_2 wl_1_2 wl_0_3
+ wl_0_4 wl_0_5 wl_1_5 wl_0_6 wl_0_7 wl_0_8 wl_1_8 wl_1_9 wl_1_10 wl_1_11 wl_1_13
+ wl_0_14 wl_1_14 wl_0_15 wl_0_16 wl_1_16 wl_0_17 wl_1_17 wl_0_18 wl_1_19 wl_1_20
+ wl_1_22 wl_1_23 wl_0_25 wl_0_26 wl_1_26 wl_0_27 wl_0_28 wl_1_28 wl_1_29 wl_1_31
+ wl_1_32 wl_1_34 wl_1_35 wl_0_36 wl_0_37 wl_1_37 wl_0_38 wl_1_38 wl_1_39 wl_1_40
+ wl_1_41 wl_1_43 wl_1_44 wl_1_46 wl_0_47 wl_1_47 wl_0_48 wl_1_49 wl_1_50 wl_1_52
+ wl_1_53 wl_0_54 wl_1_54 wl_1_55 wl_1_57 wl_0_58 wl_1_58 wl_0_59 wl_1_59 wl_1_60
+ wl_1_61 wl_0_62 wl_1_62 wl_1_63 rbl_wl_1_1 wl_0_35 wl_0_29 wl_0_20 wl_0_11 wl_0_50
+ wl_0_41 wl_0_32 wl_0_23 wl_0_53 wl_0_44 wl_1_7 rbl_wl_1_0 wl_0_46 wl_0_19 wl_0_10
+ wl_1_4 wl_0_55 wl_0_40 wl_0_31 wl_0_13 rbl_wl_0_0 wl_0_22 wl_0_57 wl_0_43 wl_0_52
+ wl_0_34 wl_1_25 wl_1_15 wl_1_6 wl_0_61 wl_0_60 wl_1_45 wl_1_36 wl_1_27 wl_1_18 wl_1_0
+ wl_0_45 wl_0_63 wl_0_9 wl_1_48 wl_1_21 wl_1_30 wl_1_12 wl_1_3 wl_0_49 wl_0_39 wl_0_30
+ wl_0_12 wl_0_21 wl_1_56 wl_1_51 wl_1_42 rbl_br_0_1 wl_1_33 wl_1_24 wl_0_56 vdd_uq0
+ wl_0_51 wl_0_42 wl_0_33 wl_0_24 rbl_bl_1_1 rbl_br_1_1 rbl_bl_0_1 gnd subbyte2_replica_column_0
.ends

.subckt subbyte2_capped_replica_bitcell_array rbl_bl_0_0 rbl_bl_1_0 rbl_br_1_0 br_1_0
+ br_1_1 br_1_2 br_1_3 bl_1_4 br_1_4 bl_1_5 br_1_5 bl_1_6 br_1_6 bl_1_7 br_1_7 bl_1_8
+ br_1_8 bl_1_9 bl_1_10 br_1_10 br_1_11 bl_1_12 br_1_12 bl_1_13 br_1_13 bl_1_14 br_1_14
+ bl_1_15 br_1_15 bl_1_16 br_1_16 bl_1_17 br_1_17 bl_1_18 br_1_18 bl_0_19 bl_1_19
+ br_0_19 bl_1_20 br_1_20 bl_1_21 br_1_21 br_1_22 bl_1_23 br_1_23 bl_1_24 br_1_24
+ bl_1_25 br_1_25 bl_1_26 br_1_26 bl_1_27 br_1_27 bl_1_28 br_1_28 bl_0_29 bl_1_29
+ bl_0_30 bl_1_30 br_1_30 bl_1_31 br_1_31 rbl_bl_0_1 rbl_bl_1_1 rbl_br_0_1 rbl_wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_1_10 wl_1_11 wl_1_12
+ wl_1_13 wl_1_14 wl_0_15 wl_1_15 wl_0_16 wl_1_16 wl_0_17 wl_1_17 wl_0_18 wl_1_18
+ wl_1_19 wl_1_20 wl_1_21 wl_1_22 wl_1_23 wl_1_24 wl_1_25 wl_0_26 wl_1_26 wl_0_27
+ wl_1_27 wl_0_28 wl_1_28 wl_1_29 wl_1_30 wl_1_31 wl_1_32 wl_1_33 wl_1_34 wl_1_35
+ wl_1_36 wl_0_37 wl_1_37 wl_0_38 wl_1_38 wl_1_39 wl_1_40 wl_1_41 wl_1_42 wl_1_43
+ wl_1_44 wl_1_45 wl_1_46 wl_1_47 wl_0_48 wl_1_48 wl_0_49 wl_1_49 wl_1_50 wl_1_51
+ wl_1_52 wl_1_53 wl_1_54 wl_1_55 wl_1_56 wl_1_57 wl_1_58 wl_0_59 wl_1_59 wl_0_60
+ wl_1_60 wl_1_61 wl_1_62 wl_1_63 rbl_wl_1_1 wl_1_9 wl_1_8 wl_1_7 wl_1_6 br_0_8 wl_1_5
+ br_0_7 br_0_18 bl_0_8 wl_1_4 br_0_6 br_0_17 br_0_28 bl_0_7 wl_1_3 br_0_5 br_0_16
+ br_0_27 bl_0_6 wl_1_2 br_0_4 br_0_15 br_0_26 bl_0_5 wl_1_1 br_0_3 br_0_25 br_0_14
+ bl_0_4 wl_1_0 br_0_2 br_0_13 br_0_24 bl_0_3 br_0_1 bl_0_18 br_0_23 br_0_12 bl_0_2
+ bl_0_17 bl_0_28 wl_0_25 wl_0_14 br_0_0 wl_0_58 wl_0_47 wl_0_36 br_0_11 br_0_22 bl_0_1
+ bl_0_16 bl_0_27 wl_0_46 wl_0_35 wl_0_13 wl_0_24 rbl_br_0_0 wl_0_57 br_0_10 br_0_21
+ bl_0_0 bl_1_3 bl_0_26 wl_0_34 wl_0_23 wl_0_56 wl_0_12 wl_0_45 bl_0_15 br_0_31 br_0_20
+ br_0_9 bl_1_2 bl_0_25 bl_0_14 wl_0_11 wl_0_55 wl_0_22 wl_0_33 wl_0_44 br_0_30 rbl_br_1_1
+ bl_1_1 bl_0_24 bl_0_13 wl_0_54 wl_0_43 wl_0_32 wl_0_21 wl_0_10 br_0_29 br_1_9 bl_1_0
+ wl_0_0 bl_0_12 bl_0_23 wl_0_31 wl_0_42 wl_0_9 wl_0_20 wl_0_53 br_1_19 bl_0_11 bl_0_22
+ wl_0_63 wl_0_30 wl_0_19 wl_0_41 wl_0_52 br_1_29 wl_0_62 wl_0_51 bl_0_10 bl_0_21
+ wl_0_29 wl_0_40 bl_0_9 wl_0_50 wl_0_39 bl_0_31 bl_0_20 wl_0_61 bl_1_11 bl_1_22 vdd
+ gnd
Xsubbyte2_replica_bitcell_array_0 bl_1_12 br_0_19 bl_1_23 wl_0_1 wl_0_2 wl_0_15 wl_0_16
+ wl_0_17 wl_0_26 wl_0_28 wl_0_37 wl_0_48 wl_0_59 vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd wl_1_44 wl_1_35 wl_1_26 br_1_24
+ bl_0_11 br_1_28 br_0_1 bl_0_22 wl_0_8 bl_0_7 bl_0_18 wl_0_35 bl_1_17 wl_0_63 wl_0_46
+ bl_1_6 wl_0_7 rbl_br_1_0 wl_0_19 bl_0_10 bl_0_21 br_0_4 wl_0_60 br_1_3 bl_1_9 br_0_25
+ wl_1_56 vdd rbl_bl_1_1 wl_1_33 wl_1_30 br_1_31 wl_1_24 wl_1_21 br_0_14 vdd rbl_wl_1_1
+ vdd vdd wl_1_15 bl_1_16 vdd wl_1_12 br_1_6 rbl_br_1_1 vdd br_1_20 bl_1_26 bl_1_15
+ wl_0_57 br_0_24 wl_0_62 wl_0_51 br_1_16 br_1_27 br_1_13 bl_0_3 br_1_12 wl_0_45 br_1_23
+ bl_1_29 bl_0_17 wl_0_13 bl_0_6 br_0_29 br_0_18 wl_0_54 bl_1_2 vdd vdd vdd wl_1_53
+ rbl_br_0_0 bl_1_0 bl_0_5 bl_1_1 gnd wl_1_50 wl_0_27 br_1_15 wl_0_10 wl_1_41 br_0_3
+ bl_0_9 br_1_26 wl_0_18 bl_1_5 bl_0_20 wl_1_47 br_0_0 br_1_2 bl_1_8 bl_0_31 bl_1_19
+ wl_0_9 bl_1_20 bl_1_4 bl_1_31 wl_0_56 wl_0_0 wl_0_42 bl_1_3 rbl_bl_0_1 br_1_29 bl_0_8
+ rbl_bl_0_0 wl_0_30 wl_0_38 br_0_31 wl_1_45 br_0_2 wl_0_24 wl_1_38 br_0_10 wl_0_21
+ wl_0_29 br_0_21 bl_0_27 wl_1_36 bl_0_23 gnd wl_1_32 wl_1_29 bl_0_16 wl_0_12 br_0_6
+ bl_0_12 rbl_br_0_1 wl_1_27 wl_1_23 bl_0_14 wl_0_6 wl_1_20 bl_0_25 bl_1_22 wl_0_3
+ br_1_5 br_0_20 bl_0_26 wl_1_18 wl_1_6 br_1_9 br_0_8 vdd wl_1_3 bl_1_11 wl_1_11 br_1_1
+ bl_1_7 br_0_9 bl_0_15 bl_1_18 wl_1_28 wl_1_9 bl_1_30 wl_1_61 wl_0_61 wl_1_58 wl_0_39
+ wl_0_52 wl_1_2 wl_0_41 br_1_0 br_0_5 wl_0_49 bl_0_30 br_0_16 wl_1_19 wl_1_0 wl_1_52
+ br_0_27 wl_1_49 wl_0_43 wl_1_57 br_0_13 wl_0_32 wl_0_40 wl_1_10 wl_1_43 br_0_12
+ wl_0_20 wl_0_55 wl_0_44 wl_0_33 wl_0_22 vdd wl_0_11 vdd wl_1_40 br_0_23 bl_0_29
+ br_1_4 wl_0_34 wl_0_23 wl_0_31 bl_1_13 br_1_22 wl_1_1 wl_1_46 wl_1_34 br_1_18 bl_1_24
+ wl_1_42 wl_1_31 bl_0_28 wl_1_39 br_1_19 bl_1_25 wl_1_55 wl_0_4 br_1_7 wl_1_17 wl_1_37
+ br_0_28 wl_1_25 br_0_11 br_0_17 br_1_17 wl_1_14 wl_0_58 wl_0_47 br_1_8 wl_0_36 bl_1_14
+ wl_0_25 wl_0_14 wl_1_22 br_0_22 wl_0_5 bl_0_2 wl_1_8 wl_1_16 wl_1_5 wl_1_13 bl_1_28
+ vdd vdd wl_1_63 bl_1_21 bl_1_10 wl_1_7 wl_0_53 bl_0_0 br_1_11 wl_1_60 bl_0_24 bl_0_13
+ wl_1_4 br_0_7 bl_0_1 br_1_10 wl_1_48 br_1_25 wl_1_54 br_0_15 br_1_21 bl_0_4 bl_1_27
+ br_0_30 bl_0_19 wl_1_62 wl_0_50 br_1_30 rbl_wl_0_0 br_0_26 wl_1_51 wl_1_59 rbl_bl_1_0
+ br_1_14 gnd subbyte2_replica_bitcell_array
.ends

.subckt subbyte2_column_mux_0 bl br bl_out br_out sel gnd
X0 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
X1 br sel br_out gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
.ends

.subckt subbyte2_column_mux_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4
+ bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12
+ br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19
+ br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26
+ br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 sel_3 bl_out_0
+ br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4
+ bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 gnd sel_2 sel_0 sel_1
Xsubbyte2_column_mux_0_0 bl_31 br_31 bl_out_7 br_out_7 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_1 bl_30 br_30 bl_out_7 br_out_7 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_2 bl_29 br_29 bl_out_7 br_out_7 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_3 bl_28 br_28 bl_out_7 br_out_7 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_4 bl_27 br_27 bl_out_6 br_out_6 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_30 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_5 bl_26 br_26 bl_out_6 br_out_6 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_20 bl_11 br_11 bl_out_2 br_out_2 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_31 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_6 bl_25 br_25 bl_out_6 br_out_6 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_10 bl_21 br_21 bl_out_5 br_out_5 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_21 bl_10 br_10 bl_out_2 br_out_2 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_7 bl_24 br_24 bl_out_6 br_out_6 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_11 bl_20 br_20 bl_out_5 br_out_5 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_22 bl_9 br_9 bl_out_2 br_out_2 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_8 bl_23 br_23 bl_out_5 br_out_5 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_12 bl_19 br_19 bl_out_4 br_out_4 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_13 bl_18 br_18 bl_out_4 br_out_4 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_23 bl_8 br_8 bl_out_2 br_out_2 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_24 bl_7 br_7 bl_out_1 br_out_1 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_9 bl_22 br_22 bl_out_5 br_out_5 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_14 bl_17 br_17 bl_out_4 br_out_4 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_25 bl_6 br_6 bl_out_1 br_out_1 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_15 bl_16 br_16 bl_out_4 br_out_4 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_26 bl_5 br_5 bl_out_1 br_out_1 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_16 bl_15 br_15 bl_out_3 br_out_3 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_27 bl_4 br_4 bl_out_1 br_out_1 sel_0 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_17 bl_14 br_14 bl_out_3 br_out_3 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_28 bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_18 bl_13 br_13 bl_out_3 br_out_3 sel_1 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_29 bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd subbyte2_column_mux_0
Xsubbyte2_column_mux_0_19 bl_12 br_12 bl_out_3 br_out_3 sel_0 gnd subbyte2_column_mux_0
.ends

.subckt sky130_fd_bd_sram__openram_sense_amp bl br dout en vdd vdd_uq0 gnd
X0 vdd_uq0 a_154_1598# dout vdd sky130_fd_pr__pfet_01v8 ad=0.3402p pd=3.06u as=0.3654p ps=3.1u w=1.26u l=0.15u
X1 a_154_1598# a_96_1989# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.8802p pd=7.6u as=0.3654p ps=3.1u w=1.26u l=0.15u
X2 gnd en a_184_1989# gnd sky130_fd_pr__nfet_01v8 ad=0.3705p pd=3.74u as=0.377p ps=3.76u w=0.65u l=0.15u
X3 a_154_1598# a_96_1989# a_184_1989# gnd sky130_fd_pr__nfet_01v8 ad=0.1885p pd=1.88u as=0p ps=0u w=0.65u l=0.15u
X4 bl en a_96_1989# vdd sky130_fd_pr__pfet_01v8 ad=0.54p pd=4.54u as=0.8802p ps=7.6u w=2u l=0.15u
X5 vdd a_154_1598# a_96_1989# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26u l=0.15u
X6 a_154_1598# en br vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0.54p ps=4.54u w=2u l=0.15u
X7 a_184_1989# a_154_1598# a_96_1989# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.1885p ps=1.88u w=0.65u l=0.15u
X8 gnd a_154_1598# dout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.1885p ps=1.88u w=0.65u l=0.15u
.ends

.subckt subbyte2_sense_amp_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4
+ data_5 bl_5 br_5 bl_6 br_6 bl_7 br_7 vdd_uq0 data_1 data_4 data_7 data_0 data_3
+ data_6 gnd vdd data_2 en
Xsky130_fd_bd_sram__openram_sense_amp_5 bl_2 br_2 data_2 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_6 bl_1 br_1 data_1 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_7 bl_0 br_0 data_0 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_1 bl_6 br_6 data_6 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_0 bl_7 br_7 data_7 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_2 bl_5 br_5 data_5 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_3 bl_4 br_4 data_4 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
Xsky130_fd_bd_sram__openram_sense_amp_4 bl_3 br_3 data_3 en vdd vdd_uq0 gnd sky130_fd_bd_sram__openram_sense_amp
.ends

.subckt subbyte2_precharge_1 bl br en_bar vdd
X0 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 ad=0.33p pd=3.4u as=0.1925p ps=1.8u w=0.55u l=0.15u
X1 vdd en_bar bl vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0.33p ps=3.4u w=0.55u l=0.15u
X2 br en_bar bl vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.55u l=0.15u
.ends

.subckt subbyte2_precharge_array_0 bl_0 br_0 bl_1 bl_3 br_3 br_4 bl_5 br_5 bl_6 br_6
+ br_7 bl_8 br_8 br_9 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 br_18 bl_19 br_19
+ br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 br_13 br_11 br_22 br_31 bl_13
+ bl_25 bl_11 bl_22 bl_31 br_1 br_23 br_12 br_20 br_32 bl_14 bl_23 bl_9 bl_12 bl_20
+ bl_32 br_2 br_10 br_24 br_21 br_30 bl_4 bl_7 bl_2 bl_10 bl_24 bl_18 bl_21 bl_30
+ en_bar vdd
Xsubbyte2_precharge_1_0 bl_32 br_32 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_1 bl_31 br_31 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_2 bl_30 br_30 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_3 bl_29 br_29 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_4 bl_28 br_28 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_5 bl_27 br_27 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_20 bl_12 br_12 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_30 bl_2 br_2 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_31 bl_1 br_1 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_6 bl_26 br_26 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_10 bl_22 br_22 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_21 bl_11 br_11 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_32 bl_0 br_0 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_7 bl_25 br_25 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_11 bl_21 br_21 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_22 bl_10 br_10 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_8 bl_24 br_24 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_12 bl_20 br_20 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_23 bl_9 br_9 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_9 bl_23 br_23 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_13 bl_19 br_19 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_24 bl_8 br_8 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_14 bl_18 br_18 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_25 bl_7 br_7 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_15 bl_17 br_17 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_26 bl_6 br_6 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_16 bl_16 br_16 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_17 bl_15 br_15 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_27 bl_5 br_5 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_28 bl_4 br_4 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_18 bl_14 br_14 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_29 bl_3 br_3 en_bar vdd subbyte2_precharge_1
Xsubbyte2_precharge_1_19 bl_13 br_13 en_bar vdd subbyte2_precharge_1
.ends

.subckt subbyte2_port_data_0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3
+ bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18
+ bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25
+ bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 dout_1 dout_2
+ dout_5 dout_6 sel_3 vdd_uq0 dout_4 sel_2 sel_1 s_en dout_0 sel_0 dout_3 vdd_uq1
+ vdd dout_7 p_en_bar gnd
Xsubbyte2_column_mux_array_0_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19
+ bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26
+ bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 sel_3 subbyte2_sense_amp_array_0/bl_0
+ subbyte2_sense_amp_array_0/br_0 subbyte2_sense_amp_array_0/bl_1 subbyte2_sense_amp_array_0/br_1
+ subbyte2_sense_amp_array_0/bl_2 subbyte2_sense_amp_array_0/br_2 subbyte2_sense_amp_array_0/bl_3
+ subbyte2_sense_amp_array_0/br_3 subbyte2_sense_amp_array_0/bl_4 subbyte2_sense_amp_array_0/br_4
+ subbyte2_sense_amp_array_0/bl_5 subbyte2_sense_amp_array_0/br_5 subbyte2_sense_amp_array_0/bl_6
+ subbyte2_sense_amp_array_0/br_6 subbyte2_sense_amp_array_0/bl_7 subbyte2_sense_amp_array_0/br_7
+ gnd sel_2 sel_0 sel_1 subbyte2_column_mux_array_0
Xsubbyte2_sense_amp_array_0 subbyte2_sense_amp_array_0/bl_0 subbyte2_sense_amp_array_0/br_0
+ subbyte2_sense_amp_array_0/bl_1 subbyte2_sense_amp_array_0/br_1 subbyte2_sense_amp_array_0/bl_2
+ subbyte2_sense_amp_array_0/br_2 subbyte2_sense_amp_array_0/bl_3 subbyte2_sense_amp_array_0/br_3
+ subbyte2_sense_amp_array_0/bl_4 subbyte2_sense_amp_array_0/br_4 dout_5 subbyte2_sense_amp_array_0/bl_5
+ subbyte2_sense_amp_array_0/br_5 subbyte2_sense_amp_array_0/bl_6 subbyte2_sense_amp_array_0/br_6
+ subbyte2_sense_amp_array_0/bl_7 subbyte2_sense_amp_array_0/br_7 vdd_uq1 dout_1 dout_4
+ dout_7 dout_0 dout_3 dout_6 gnd vdd dout_2 s_en subbyte2_sense_amp_array
Xsubbyte2_precharge_array_0_0 bl_0 br_0 bl_1 bl_3 br_3 br_4 bl_5 br_5 bl_6 br_6 br_7
+ bl_8 br_8 br_9 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 br_18 bl_19 br_19 br_25
+ bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 br_13 br_11 br_22 br_31 bl_13 bl_25
+ bl_11 bl_22 bl_31 br_1 br_23 br_12 br_20 rbl_br bl_14 bl_23 bl_9 bl_12 bl_20 rbl_bl
+ br_2 br_10 br_24 br_21 br_30 bl_4 bl_7 bl_2 bl_10 bl_24 bl_18 bl_21 bl_30 p_en_bar
+ vdd_uq0 subbyte2_precharge_array_0
.ends

.subckt subbyte2_precharge_0 bl br en_bar vdd
X0 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 ad=0.33p pd=3.4u as=0.1925p ps=1.8u w=0.55u l=0.15u
X1 vdd en_bar bl vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0.33p ps=3.4u w=0.55u l=0.15u
X2 br en_bar bl vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.55u l=0.15u
.ends

.subckt subbyte2_precharge_array bl_0 bl_1 bl_3 br_3 br_4 bl_5 bl_6 br_6 br_7 bl_8
+ br_8 bl_9 br_9 br_11 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19
+ br_19 br_25 bl_26 br_26 bl_27 br_27 br_28 bl_29 br_29 br_13 br_22 br_23 br_32 bl_13
+ bl_11 bl_22 bl_23 bl_32 br_1 br_12 br_20 br_24 br_30 bl_14 bl_12 bl_20 bl_24 bl_30
+ br_2 br_10 br_21 br_31 bl_4 bl_7 bl_2 bl_10 bl_21 bl_25 vdd bl_28 bl_31 br_0 br_5
+ en_bar
Xsubbyte2_precharge_0_13 bl_19 br_19 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_24 bl_8 br_8 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_14 bl_18 br_18 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_25 bl_7 br_7 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_15 bl_17 br_17 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_26 bl_6 br_6 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_16 bl_16 br_16 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_27 bl_5 br_5 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_17 bl_15 br_15 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_28 bl_4 br_4 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_18 bl_14 br_14 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_19 bl_13 br_13 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_29 bl_3 br_3 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_0 bl_32 br_32 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_1 bl_31 br_31 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_2 bl_30 br_30 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_3 bl_29 br_29 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_4 bl_28 br_28 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_5 bl_27 br_27 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_6 bl_26 br_26 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_7 bl_25 br_25 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_8 bl_24 br_24 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_9 bl_23 br_23 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_30 bl_2 br_2 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_10 bl_22 br_22 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_20 bl_12 br_12 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_21 bl_11 br_11 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_31 bl_1 br_1 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_32 bl_0 br_0 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_11 bl_21 br_21 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_22 bl_10 br_10 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_12 bl_20 br_20 en_bar vdd subbyte2_precharge_0
Xsubbyte2_precharge_0_23 bl_9 br_9 en_bar vdd subbyte2_precharge_0
.ends

.subckt sky130_fd_bd_sram__openram_write_driver din bl br en vdd gnd vdd_uq0
X0 a_213_736# en a_129_736# gnd sky130_fd_pr__nfet_01v8 ad=0.1595p pd=1.68u as=0.1485p ps=1.64u w=0.55u l=0.15u
X1 a_271_690# din gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1044p pd=1.3u as=0.7312p ps=7.36u w=0.36u l=0.15u
X2 vdd a_41_1120# a_121_1585# vdd sky130_fd_pr__pfet_01v8 ad=0.319p pd=3.36u as=0.1485p ps=1.64u w=0.55u l=0.15u
X3 a_271_690# din vdd_uq0 vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0.15125p pd=1.65u as=0.308p ps=3.32u w=0.55u l=0.15u
X4 a_129_736# a_271_690# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29975p pd=3.29u as=0p ps=0u w=0.55u l=0.15u
X5 a_41_1120# en vdd_uq0 vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0.1595p pd=1.68u as=0p ps=0u w=0.55u l=0.15u
X6 br a_121_1585# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.27p pd=2.54u as=0p ps=0u w=1u l=0.15u
X7 a_183_1687# a_129_736# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0972p pd=1.26u as=0p ps=0u w=0.36u l=0.15u
X8 gnd din a_145_492# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.1595p ps=1.68u w=0.55u l=0.15u
X9 vdd en a_129_736# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.55u l=0.15u
X10 gnd a_271_690# a_213_736# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.55u l=0.15u
X11 a_183_1687# a_129_736# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1485p pd=1.64u as=0p ps=0u w=0.55u l=0.15u
X12 gnd a_183_1687# bl gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.27p ps=2.54u w=1u l=0.15u
X13 gnd a_41_1120# a_121_1585# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.0972p ps=1.26u w=0.36u l=0.15u
X14 vdd_uq0 din a_41_1120# vdd_uq0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.55u l=0.15u
X15 a_145_492# en a_41_1120# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0.1485p ps=1.64u w=0.55u l=0.15u
.ends

.subckt subbyte2_write_driver_array data_1 data_4 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3
+ br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 vdd_uq0 data_7 data_0 data_3 data_6
+ data_2 data_5 gnd en vdd
Xsky130_fd_bd_sram__openram_write_driver_7 data_0 bl_0 br_0 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_0 data_7 bl_7 br_7 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_1 data_6 bl_6 br_6 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_2 data_5 bl_5 br_5 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_3 data_4 bl_4 br_4 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_5 data_2 bl_2 br_2 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_4 data_3 bl_3 br_3 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
Xsky130_fd_bd_sram__openram_write_driver_6 data_1 bl_1 br_1 en vdd gnd vdd_uq0 sky130_fd_bd_sram__openram_write_driver
.ends

.subckt subbyte2_column_mux bl br bl_out br_out sel gnd
X0 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
X1 br sel br_out gnd sky130_fd_pr__nfet_01v8 ad=0.864p pd=6.36u as=0.864p ps=6.36u w=2.88u l=0.15u
.ends

.subckt subbyte2_column_mux_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4
+ bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12
+ br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19
+ br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26
+ br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 sel_3 bl_out_0
+ br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4
+ bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 sel_2 sel_1 gnd sel_0
Xsubbyte2_column_mux_30 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_20 bl_11 br_11 bl_out_2 br_out_2 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_31 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_10 bl_21 br_21 bl_out_5 br_out_5 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_21 bl_10 br_10 bl_out_2 br_out_2 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_11 bl_20 br_20 bl_out_5 br_out_5 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_22 bl_9 br_9 bl_out_2 br_out_2 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_12 bl_19 br_19 bl_out_4 br_out_4 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_23 bl_8 br_8 bl_out_2 br_out_2 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_13 bl_18 br_18 bl_out_4 br_out_4 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_24 bl_7 br_7 bl_out_1 br_out_1 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_14 bl_17 br_17 bl_out_4 br_out_4 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_25 bl_6 br_6 bl_out_1 br_out_1 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_15 bl_16 br_16 bl_out_4 br_out_4 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_26 bl_5 br_5 bl_out_1 br_out_1 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_16 bl_15 br_15 bl_out_3 br_out_3 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_17 bl_14 br_14 bl_out_3 br_out_3 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_27 bl_4 br_4 bl_out_1 br_out_1 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_28 bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_18 bl_13 br_13 bl_out_3 br_out_3 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_29 bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_0 bl_31 br_31 bl_out_7 br_out_7 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_19 bl_12 br_12 bl_out_3 br_out_3 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_1 bl_30 br_30 bl_out_7 br_out_7 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_2 bl_29 br_29 bl_out_7 br_out_7 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_3 bl_28 br_28 bl_out_7 br_out_7 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_4 bl_27 br_27 bl_out_6 br_out_6 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_5 bl_26 br_26 bl_out_6 br_out_6 sel_2 gnd subbyte2_column_mux
Xsubbyte2_column_mux_6 bl_25 br_25 bl_out_6 br_out_6 sel_1 gnd subbyte2_column_mux
Xsubbyte2_column_mux_7 bl_24 br_24 bl_out_6 br_out_6 sel_0 gnd subbyte2_column_mux
Xsubbyte2_column_mux_8 bl_23 br_23 bl_out_5 br_out_5 sel_3 gnd subbyte2_column_mux
Xsubbyte2_column_mux_9 bl_22 br_22 bl_out_5 br_out_5 sel_2 gnd subbyte2_column_mux
.ends

.subckt subbyte2_port_data rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4
+ br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12
+ br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19
+ br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26
+ br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 din_7 sel_3 din_2
+ din_1 din_4 din_5 sel_2 sel_1 sel_0 w_en din_0 din_3 p_en_bar vdd din_6 vdd_uq1
+ vdd_uq0 gnd
Xsubbyte2_precharge_array_0 rbl_bl bl_0 bl_2 br_2 br_3 bl_4 bl_5 br_5 br_6 bl_7 br_7
+ bl_8 br_8 br_10 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18
+ br_24 bl_25 br_25 bl_26 br_26 br_27 bl_28 br_28 br_12 br_21 br_22 br_31 bl_12 bl_10
+ bl_21 bl_22 bl_31 br_0 br_11 br_19 br_23 br_29 bl_13 bl_11 bl_19 bl_23 bl_29 br_1
+ br_9 br_20 br_30 bl_3 bl_6 bl_1 bl_9 bl_20 bl_24 vdd_uq0 bl_27 bl_30 rbl_br br_4
+ p_en_bar subbyte2_precharge_array
Xsubbyte2_write_driver_array_0 din_1 din_4 subbyte2_write_driver_array_0/bl_0 subbyte2_write_driver_array_0/br_0
+ subbyte2_write_driver_array_0/bl_1 subbyte2_write_driver_array_0/br_1 subbyte2_write_driver_array_0/bl_2
+ subbyte2_write_driver_array_0/br_2 subbyte2_write_driver_array_0/bl_3 subbyte2_write_driver_array_0/br_3
+ subbyte2_write_driver_array_0/bl_4 subbyte2_write_driver_array_0/br_4 subbyte2_write_driver_array_0/bl_5
+ subbyte2_write_driver_array_0/br_5 subbyte2_write_driver_array_0/bl_6 subbyte2_write_driver_array_0/br_6
+ subbyte2_write_driver_array_0/bl_7 subbyte2_write_driver_array_0/br_7 vdd_uq1 din_7
+ din_0 din_3 din_6 din_2 din_5 gnd w_en vdd subbyte2_write_driver_array
Xsubbyte2_column_mux_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19
+ bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26
+ bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 sel_3 subbyte2_write_driver_array_0/bl_0
+ subbyte2_write_driver_array_0/br_0 subbyte2_write_driver_array_0/bl_1 subbyte2_write_driver_array_0/br_1
+ subbyte2_write_driver_array_0/bl_2 subbyte2_write_driver_array_0/br_2 subbyte2_write_driver_array_0/bl_3
+ subbyte2_write_driver_array_0/br_3 subbyte2_write_driver_array_0/bl_4 subbyte2_write_driver_array_0/br_4
+ subbyte2_write_driver_array_0/bl_5 subbyte2_write_driver_array_0/br_5 subbyte2_write_driver_array_0/bl_6
+ subbyte2_write_driver_array_0/br_6 subbyte2_write_driver_array_0/bl_7 subbyte2_write_driver_array_0/br_7
+ sel_2 sel_1 gnd sel_0 subbyte2_column_mux_array
.ends

.subckt subbyte2_pinv_dec_0 A Z vdd gnd
X0 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.9p pd=6.6u as=0.9p ps=6.6u w=3u l=0.15u
X1 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=2.1p pd=14.6u as=2.1p ps=14.6u w=7u l=0.15u
.ends

.subckt sky130_fd_bd_sram__openram_dp_nand2_dec A B Z gnd vdd
X0 Z A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.6048p pd=5.56u as=0.336p ps=2.84u w=1.12u l=0.15u
X1 vdd B Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X2 a_196_224# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1554p pd=1.9u as=0.3182p ps=2.34u w=0.74u l=0.15u
X3 Z A a_196_224# gnd sky130_fd_pr__nfet_01v8 ad=0.222p pd=2.08u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt subbyte2_and2_dec_0 A B Z vdd_uq0 vdd gnd
Xsubbyte2_pinv_dec_0_0 subbyte2_pinv_dec_0_0/A Z vdd_uq0 gnd subbyte2_pinv_dec_0
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B subbyte2_pinv_dec_0_0/A gnd vdd sky130_fd_bd_sram__openram_dp_nand2_dec
.ends

.subckt sky130_fd_bd_sram__openram_dp_nand3_dec A B C Z gnd vdd
X0 Z B vdd vdd sky130_fd_pr__pfet_01v8 ad=1.008p pd=8.52u as=0.7728p ps=5.86u w=1.12u l=0.15u
X1 vdd C Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X2 a_198_136# A Z gnd sky130_fd_pr__nfet_01v8 ad=0.1554p pd=1.9u as=0.222p ps=2.08u w=0.74u l=0.15u
X3 gnd C a_198_208# gnd sky130_fd_pr__nfet_01v8 ad=0.3108p pd=2.32u as=0.1554p ps=1.9u w=0.74u l=0.15u
X4 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12u l=0.15u
X5 a_198_208# B a_198_136# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0.74u l=0.15u
.ends

.subckt subbyte2_pinv_dec A Z vdd gnd
X0 gnd A Z gnd sky130_fd_pr__nfet_01v8 ad=0.108p pd=1.32u as=0.108p ps=1.32u w=0.36u l=0.15u
X1 vdd A Z vdd sky130_fd_pr__pfet_01v8 ad=0.336p pd=2.84u as=0.336p ps=2.84u w=1.12u l=0.15u
.ends

.subckt subbyte2_and3_dec A vdd_uq0 vdd gnd C B Z
Xsky130_fd_bd_sram__openram_dp_nand3_dec_0 A B C subbyte2_pinv_dec_0/A gnd vdd sky130_fd_bd_sram__openram_dp_nand3_dec
Xsubbyte2_pinv_dec_0 subbyte2_pinv_dec_0/A Z vdd_uq0 gnd subbyte2_pinv_dec
.ends

.subckt subbyte2_and2_dec A B Z vdd_uq0 vdd gnd
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B subbyte2_pinv_dec_0/A gnd vdd sky130_fd_bd_sram__openram_dp_nand2_dec
Xsubbyte2_pinv_dec_0 subbyte2_pinv_dec_0/A Z vdd_uq0 gnd subbyte2_pinv_dec
.ends

.subckt subbyte2_hierarchical_predecode2x4 in_0 in_1 out_0 out_1 out_2 out_3 vdd_uq0
+ vdd_uq1 gnd vdd
Xsubbyte2_and2_dec_0 in_0 in_1 out_3 vdd_uq0 vdd gnd subbyte2_and2_dec
Xsubbyte2_and2_dec_2 in_0 subbyte2_pinv_dec_0/Z out_1 vdd_uq0 vdd gnd subbyte2_and2_dec
Xsubbyte2_and2_dec_1 subbyte2_pinv_dec_1/Z in_1 out_2 vdd_uq0 vdd gnd subbyte2_and2_dec
Xsubbyte2_and2_dec_3 subbyte2_pinv_dec_1/Z subbyte2_pinv_dec_0/Z out_0 vdd_uq0 vdd
+ gnd subbyte2_and2_dec
Xsubbyte2_pinv_dec_0 in_1 subbyte2_pinv_dec_0/Z vdd_uq1 gnd subbyte2_pinv_dec
Xsubbyte2_pinv_dec_1 in_0 subbyte2_pinv_dec_1/Z vdd_uq1 gnd subbyte2_pinv_dec
.ends

.subckt subbyte2_hierarchical_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 decode_0
+ decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9
+ decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17
+ decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25
+ decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33
+ decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41
+ decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49
+ decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57
+ decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 vdd_uq2 vdd_uq1 vdd
+ vdd_uq7 vdd_uq8 vdd_uq6 vdd_uq9 vdd_uq11 vdd_uq13 vdd_uq14 vdd_uq16 gnd
Xsubbyte2_and3_dec_12 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_63/B decode_51 subbyte2_and3_dec
Xsubbyte2_and3_dec_23 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_7/B decode_40 subbyte2_and3_dec
Xsubbyte2_and3_dec_34 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_3/B decode_29 subbyte2_and3_dec
Xsubbyte2_and3_dec_45 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_63/B decode_18 subbyte2_and3_dec
Xsubbyte2_and3_dec_56 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_9/B decode_7 subbyte2_and3_dec
Xsubbyte2_and3_dec_13 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_63/B decode_50 subbyte2_and3_dec
Xsubbyte2_and3_dec_24 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_9/B decode_39 subbyte2_and3_dec
Xsubbyte2_and3_dec_35 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_3/B decode_28 subbyte2_and3_dec
Xsubbyte2_and3_dec_46 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_63/B decode_17 subbyte2_and3_dec
Xsubbyte2_and3_dec_57 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_9/B decode_6 subbyte2_and3_dec
Xsubbyte2_and3_dec_14 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_63/B decode_49 subbyte2_and3_dec
Xsubbyte2_and3_dec_25 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_9/B decode_38 subbyte2_and3_dec
Xsubbyte2_and3_dec_36 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_7/B decode_27 subbyte2_and3_dec
Xsubbyte2_and3_dec_47 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_63/B decode_16 subbyte2_and3_dec
Xsubbyte2_and3_dec_58 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_9/B decode_5 subbyte2_and3_dec
Xsubbyte2_and3_dec_15 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_63/B decode_48 subbyte2_and3_dec
Xsubbyte2_and3_dec_26 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_9/B decode_37 subbyte2_and3_dec
Xsubbyte2_and3_dec_37 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_7/B decode_26 subbyte2_and3_dec
Xsubbyte2_and3_dec_48 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_3/B decode_15 subbyte2_and3_dec
Xsubbyte2_and3_dec_59 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_9/B decode_4 subbyte2_and3_dec
Xsubbyte2_and3_dec_16 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_3/B decode_47 subbyte2_and3_dec
Xsubbyte2_and3_dec_27 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_9/B decode_36 subbyte2_and3_dec
Xsubbyte2_and3_dec_38 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_7/B decode_25 subbyte2_and3_dec
Xsubbyte2_and3_dec_49 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_3/B decode_14 subbyte2_and3_dec
Xsubbyte2_and3_dec_17 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_3/B decode_46 subbyte2_and3_dec
Xsubbyte2_and3_dec_28 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_63/B decode_35 subbyte2_and3_dec
Xsubbyte2_and3_dec_39 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_7/B decode_24 subbyte2_and3_dec
Xsubbyte2_and3_dec_18 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_3/B decode_45 subbyte2_and3_dec
Xsubbyte2_and3_dec_19 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_3/B decode_44 subbyte2_and3_dec
Xsubbyte2_and3_dec_29 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_63/B decode_34 subbyte2_and3_dec
Xsubbyte2_hierarchical_predecode2x4_0 addr_4 addr_5 subbyte2_and3_dec_63/C subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_31/C subbyte2_and3_dec_9/C vdd_uq9 vdd_uq11 gnd vdd_uq13 subbyte2_hierarchical_predecode2x4
Xsubbyte2_hierarchical_predecode2x4_1 addr_2 addr_3 subbyte2_and3_dec_63/B subbyte2_and3_dec_9/B
+ subbyte2_and3_dec_7/B subbyte2_and3_dec_3/B vdd_uq7 vdd_uq6 gnd vdd_uq8 subbyte2_hierarchical_predecode2x4
Xsubbyte2_hierarchical_predecode2x4_2 addr_0 addr_1 subbyte2_and3_dec_7/A subbyte2_and3_dec_6/A
+ subbyte2_and3_dec_9/A subbyte2_and3_dec_8/A vdd_uq2 vdd_uq1 gnd vdd subbyte2_hierarchical_predecode2x4
Xsubbyte2_and3_dec_0 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_3/B decode_63 subbyte2_and3_dec
Xsubbyte2_and3_dec_1 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_3/B decode_62 subbyte2_and3_dec
Xsubbyte2_and3_dec_2 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_3/B decode_61 subbyte2_and3_dec
Xsubbyte2_and3_dec_3 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_3/B decode_60 subbyte2_and3_dec
Xsubbyte2_and3_dec_4 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_7/B decode_59 subbyte2_and3_dec
Xsubbyte2_and3_dec_5 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_7/B decode_58 subbyte2_and3_dec
Xsubbyte2_and3_dec_6 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_7/B decode_57 subbyte2_and3_dec
Xsubbyte2_and3_dec_7 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_7/B decode_56 subbyte2_and3_dec
Xsubbyte2_and3_dec_60 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_63/B decode_3 subbyte2_and3_dec
Xsubbyte2_and3_dec_8 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_9/B decode_55 subbyte2_and3_dec
Xsubbyte2_and3_dec_50 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_3/B decode_13 subbyte2_and3_dec
Xsubbyte2_and3_dec_61 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_63/B decode_2 subbyte2_and3_dec
Xsubbyte2_and3_dec_9 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_9/B decode_54 subbyte2_and3_dec
Xsubbyte2_and3_dec_40 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_9/B decode_23 subbyte2_and3_dec
Xsubbyte2_and3_dec_51 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_3/B decode_12 subbyte2_and3_dec
Xsubbyte2_and3_dec_62 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_63/B decode_1 subbyte2_and3_dec
Xsubbyte2_and3_dec_30 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_63/B decode_33 subbyte2_and3_dec
Xsubbyte2_and3_dec_41 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_9/B decode_22 subbyte2_and3_dec
Xsubbyte2_and3_dec_52 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_7/B decode_11 subbyte2_and3_dec
Xsubbyte2_and3_dec_63 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_63/B decode_0 subbyte2_and3_dec
Xsubbyte2_and3_dec_10 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_9/B decode_53 subbyte2_and3_dec
Xsubbyte2_and3_dec_20 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_7/B decode_43 subbyte2_and3_dec
Xsubbyte2_and3_dec_21 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_7/B decode_42 subbyte2_and3_dec
Xsubbyte2_and3_dec_31 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_63/B decode_32 subbyte2_and3_dec
Xsubbyte2_and3_dec_32 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_3/B decode_31 subbyte2_and3_dec
Xsubbyte2_and3_dec_42 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_9/B decode_21 subbyte2_and3_dec
Xsubbyte2_and3_dec_43 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_9/B decode_20 subbyte2_and3_dec
Xsubbyte2_and3_dec_53 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_7/B decode_10 subbyte2_and3_dec
Xsubbyte2_and3_dec_54 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_7/B decode_9 subbyte2_and3_dec
Xsubbyte2_and3_dec_11 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_9/C
+ subbyte2_and3_dec_9/B decode_52 subbyte2_and3_dec
Xsubbyte2_and3_dec_22 subbyte2_and3_dec_6/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_31/C
+ subbyte2_and3_dec_7/B decode_41 subbyte2_and3_dec
Xsubbyte2_and3_dec_33 subbyte2_and3_dec_9/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_3/B decode_30 subbyte2_and3_dec
Xsubbyte2_and3_dec_44 subbyte2_and3_dec_8/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_47/C
+ subbyte2_and3_dec_63/B decode_19 subbyte2_and3_dec
Xsubbyte2_and3_dec_55 subbyte2_and3_dec_7/A vdd_uq14 vdd_uq16 gnd subbyte2_and3_dec_63/C
+ subbyte2_and3_dec_7/B decode_8 subbyte2_and3_dec
.ends

.subckt subbyte2_wordline_driver Z vdd_uq0 B A vdd gnd
Xsubbyte2_pinv_dec_0_0 subbyte2_pinv_dec_0_0/A Z vdd_uq0 gnd subbyte2_pinv_dec_0
Xsky130_fd_bd_sram__openram_dp_nand2_dec_0 A B subbyte2_pinv_dec_0_0/A gnd vdd sky130_fd_bd_sram__openram_dp_nand2_dec
.ends

.subckt subbyte2_wordline_driver_array in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8
+ in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22
+ in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36
+ in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50
+ in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43
+ wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57
+ wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 en vdd vdd_uq0 gnd
Xsubbyte2_wordline_driver_7 wl_56 vdd_uq0 en in_56 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_8 wl_55 vdd_uq0 en in_55 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_9 wl_54 vdd_uq0 en in_54 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_60 wl_3 vdd_uq0 en in_3 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_50 wl_13 vdd_uq0 en in_13 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_61 wl_2 vdd_uq0 en in_2 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_40 wl_23 vdd_uq0 en in_23 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_51 wl_12 vdd_uq0 en in_12 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_62 wl_1 vdd_uq0 en in_1 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_30 wl_33 vdd_uq0 en in_33 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_41 wl_22 vdd_uq0 en in_22 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_52 wl_11 vdd_uq0 en in_11 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_63 wl_0 vdd_uq0 en in_0 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_20 wl_43 vdd_uq0 en in_43 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_31 wl_32 vdd_uq0 en in_32 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_42 wl_21 vdd_uq0 en in_21 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_53 wl_10 vdd_uq0 en in_10 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_10 wl_53 vdd_uq0 en in_53 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_21 wl_42 vdd_uq0 en in_42 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_32 wl_31 vdd_uq0 en in_31 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_43 wl_20 vdd_uq0 en in_20 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_54 wl_9 vdd_uq0 en in_9 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_11 wl_52 vdd_uq0 en in_52 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_12 wl_51 vdd_uq0 en in_51 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_22 wl_41 vdd_uq0 en in_41 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_23 wl_40 vdd_uq0 en in_40 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_33 wl_30 vdd_uq0 en in_30 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_34 wl_29 vdd_uq0 en in_29 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_44 wl_19 vdd_uq0 en in_19 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_55 wl_8 vdd_uq0 en in_8 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_13 wl_50 vdd_uq0 en in_50 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_24 wl_39 vdd_uq0 en in_39 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_35 wl_28 vdd_uq0 en in_28 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_45 wl_18 vdd_uq0 en in_18 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_46 wl_17 vdd_uq0 en in_17 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_56 wl_7 vdd_uq0 en in_7 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_57 wl_6 vdd_uq0 en in_6 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_14 wl_49 vdd_uq0 en in_49 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_25 wl_38 vdd_uq0 en in_38 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_36 wl_27 vdd_uq0 en in_27 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_47 wl_16 vdd_uq0 en in_16 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_58 wl_5 vdd_uq0 en in_5 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_15 wl_48 vdd_uq0 en in_48 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_26 wl_37 vdd_uq0 en in_37 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_37 wl_26 vdd_uq0 en in_26 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_48 wl_15 vdd_uq0 en in_15 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_59 wl_4 vdd_uq0 en in_4 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_16 wl_47 vdd_uq0 en in_47 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_27 wl_36 vdd_uq0 en in_36 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_38 wl_25 vdd_uq0 en in_25 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_49 wl_14 vdd_uq0 en in_14 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_17 wl_46 vdd_uq0 en in_46 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_28 wl_35 vdd_uq0 en in_35 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_39 wl_24 vdd_uq0 en in_24 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_18 wl_45 vdd_uq0 en in_45 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_29 wl_34 vdd_uq0 en in_34 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_19 wl_44 vdd_uq0 en in_44 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_0 wl_63 vdd_uq0 en in_63 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_1 wl_62 vdd_uq0 en in_62 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_2 wl_61 vdd_uq0 en in_61 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_3 wl_60 vdd_uq0 en in_60 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_4 wl_59 vdd_uq0 en in_59 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_5 wl_58 vdd_uq0 en in_58 vdd gnd subbyte2_wordline_driver
Xsubbyte2_wordline_driver_6 wl_57 vdd_uq0 en in_57 vdd gnd subbyte2_wordline_driver
.ends

.subckt subbyte2_port_address addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 wl_en wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43
+ wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57
+ wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 rbl_wl vdd_uq7 vdd_uq8 vdd_uq6 vdd_uq21 vdd_uq17
+ vdd_uq16 vdd_uq11 vdd_uq9 vdd_uq13 vdd_uq18 vdd_uq0 vdd vdd_uq3 vdd_uq1 gnd
Xsubbyte2_and2_dec_0_0 wl_en vdd_uq21 rbl_wl vdd_uq0 vdd gnd subbyte2_and2_dec_0
Xsubbyte2_hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 subbyte2_wordline_driver_array_0/in_0
+ subbyte2_wordline_driver_array_0/in_1 subbyte2_wordline_driver_array_0/in_2 subbyte2_wordline_driver_array_0/in_3
+ subbyte2_wordline_driver_array_0/in_4 subbyte2_wordline_driver_array_0/in_5 subbyte2_wordline_driver_array_0/in_6
+ subbyte2_wordline_driver_array_0/in_7 subbyte2_wordline_driver_array_0/in_8 subbyte2_wordline_driver_array_0/in_9
+ subbyte2_wordline_driver_array_0/in_10 subbyte2_wordline_driver_array_0/in_11 subbyte2_wordline_driver_array_0/in_12
+ subbyte2_wordline_driver_array_0/in_13 subbyte2_wordline_driver_array_0/in_14 subbyte2_wordline_driver_array_0/in_15
+ subbyte2_wordline_driver_array_0/in_16 subbyte2_wordline_driver_array_0/in_17 subbyte2_wordline_driver_array_0/in_18
+ subbyte2_wordline_driver_array_0/in_19 subbyte2_wordline_driver_array_0/in_20 subbyte2_wordline_driver_array_0/in_21
+ subbyte2_wordline_driver_array_0/in_22 subbyte2_wordline_driver_array_0/in_23 subbyte2_wordline_driver_array_0/in_24
+ subbyte2_wordline_driver_array_0/in_25 subbyte2_wordline_driver_array_0/in_26 subbyte2_wordline_driver_array_0/in_27
+ subbyte2_wordline_driver_array_0/in_28 subbyte2_wordline_driver_array_0/in_29 subbyte2_wordline_driver_array_0/in_30
+ subbyte2_wordline_driver_array_0/in_31 subbyte2_wordline_driver_array_0/in_32 subbyte2_wordline_driver_array_0/in_33
+ subbyte2_wordline_driver_array_0/in_34 subbyte2_wordline_driver_array_0/in_35 subbyte2_wordline_driver_array_0/in_36
+ subbyte2_wordline_driver_array_0/in_37 subbyte2_wordline_driver_array_0/in_38 subbyte2_wordline_driver_array_0/in_39
+ subbyte2_wordline_driver_array_0/in_40 subbyte2_wordline_driver_array_0/in_41 subbyte2_wordline_driver_array_0/in_42
+ subbyte2_wordline_driver_array_0/in_43 subbyte2_wordline_driver_array_0/in_44 subbyte2_wordline_driver_array_0/in_45
+ subbyte2_wordline_driver_array_0/in_46 subbyte2_wordline_driver_array_0/in_47 subbyte2_wordline_driver_array_0/in_48
+ subbyte2_wordline_driver_array_0/in_49 subbyte2_wordline_driver_array_0/in_50 subbyte2_wordline_driver_array_0/in_51
+ subbyte2_wordline_driver_array_0/in_52 subbyte2_wordline_driver_array_0/in_53 subbyte2_wordline_driver_array_0/in_54
+ subbyte2_wordline_driver_array_0/in_55 subbyte2_wordline_driver_array_0/in_56 subbyte2_wordline_driver_array_0/in_57
+ subbyte2_wordline_driver_array_0/in_58 subbyte2_wordline_driver_array_0/in_59 subbyte2_wordline_driver_array_0/in_60
+ subbyte2_wordline_driver_array_0/in_61 subbyte2_wordline_driver_array_0/in_62 subbyte2_wordline_driver_array_0/in_63
+ vdd_uq7 vdd_uq6 vdd_uq8 vdd_uq9 vdd_uq13 vdd_uq11 vdd_uq17 vdd_uq16 vdd_uq18 vdd_uq1
+ vdd_uq3 gnd subbyte2_hierarchical_decoder
Xsubbyte2_wordline_driver_array_0 subbyte2_wordline_driver_array_0/in_0 subbyte2_wordline_driver_array_0/in_1
+ subbyte2_wordline_driver_array_0/in_2 subbyte2_wordline_driver_array_0/in_3 subbyte2_wordline_driver_array_0/in_4
+ subbyte2_wordline_driver_array_0/in_5 subbyte2_wordline_driver_array_0/in_6 subbyte2_wordline_driver_array_0/in_7
+ subbyte2_wordline_driver_array_0/in_8 subbyte2_wordline_driver_array_0/in_9 subbyte2_wordline_driver_array_0/in_10
+ subbyte2_wordline_driver_array_0/in_11 subbyte2_wordline_driver_array_0/in_12 subbyte2_wordline_driver_array_0/in_13
+ subbyte2_wordline_driver_array_0/in_14 subbyte2_wordline_driver_array_0/in_15 subbyte2_wordline_driver_array_0/in_16
+ subbyte2_wordline_driver_array_0/in_17 subbyte2_wordline_driver_array_0/in_18 subbyte2_wordline_driver_array_0/in_19
+ subbyte2_wordline_driver_array_0/in_20 subbyte2_wordline_driver_array_0/in_21 subbyte2_wordline_driver_array_0/in_22
+ subbyte2_wordline_driver_array_0/in_23 subbyte2_wordline_driver_array_0/in_24 subbyte2_wordline_driver_array_0/in_25
+ subbyte2_wordline_driver_array_0/in_26 subbyte2_wordline_driver_array_0/in_27 subbyte2_wordline_driver_array_0/in_28
+ subbyte2_wordline_driver_array_0/in_29 subbyte2_wordline_driver_array_0/in_30 subbyte2_wordline_driver_array_0/in_31
+ subbyte2_wordline_driver_array_0/in_32 subbyte2_wordline_driver_array_0/in_33 subbyte2_wordline_driver_array_0/in_34
+ subbyte2_wordline_driver_array_0/in_35 subbyte2_wordline_driver_array_0/in_36 subbyte2_wordline_driver_array_0/in_37
+ subbyte2_wordline_driver_array_0/in_38 subbyte2_wordline_driver_array_0/in_39 subbyte2_wordline_driver_array_0/in_40
+ subbyte2_wordline_driver_array_0/in_41 subbyte2_wordline_driver_array_0/in_42 subbyte2_wordline_driver_array_0/in_43
+ subbyte2_wordline_driver_array_0/in_44 subbyte2_wordline_driver_array_0/in_45 subbyte2_wordline_driver_array_0/in_46
+ subbyte2_wordline_driver_array_0/in_47 subbyte2_wordline_driver_array_0/in_48 subbyte2_wordline_driver_array_0/in_49
+ subbyte2_wordline_driver_array_0/in_50 subbyte2_wordline_driver_array_0/in_51 subbyte2_wordline_driver_array_0/in_52
+ subbyte2_wordline_driver_array_0/in_53 subbyte2_wordline_driver_array_0/in_54 subbyte2_wordline_driver_array_0/in_55
+ subbyte2_wordline_driver_array_0/in_56 subbyte2_wordline_driver_array_0/in_57 subbyte2_wordline_driver_array_0/in_58
+ subbyte2_wordline_driver_array_0/in_59 subbyte2_wordline_driver_array_0/in_60 subbyte2_wordline_driver_array_0/in_61
+ subbyte2_wordline_driver_array_0/in_62 subbyte2_wordline_driver_array_0/in_63 wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43
+ wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57
+ wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_en vdd vdd_uq0 gnd subbyte2_wordline_driver_array
.ends

.subckt subbyte2_port_address_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 wl_en wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43
+ wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57
+ wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 rbl_wl vdd_uq3 vdd_uq7 vdd_uq8 vdd_uq6 vdd_uq21
+ vdd_uq17 vdd_uq16 vdd_uq11 vdd_uq9 vdd_uq13 vdd_uq18 vdd_uq0 vdd gnd vdd_uq1
Xsubbyte2_and2_dec_0_0 wl_en vdd_uq21 rbl_wl vdd_uq0 vdd gnd subbyte2_and2_dec_0
Xsubbyte2_hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 subbyte2_wordline_driver_array_0/in_0
+ subbyte2_wordline_driver_array_0/in_1 subbyte2_wordline_driver_array_0/in_2 subbyte2_wordline_driver_array_0/in_3
+ subbyte2_wordline_driver_array_0/in_4 subbyte2_wordline_driver_array_0/in_5 subbyte2_wordline_driver_array_0/in_6
+ subbyte2_wordline_driver_array_0/in_7 subbyte2_wordline_driver_array_0/in_8 subbyte2_wordline_driver_array_0/in_9
+ subbyte2_wordline_driver_array_0/in_10 subbyte2_wordline_driver_array_0/in_11 subbyte2_wordline_driver_array_0/in_12
+ subbyte2_wordline_driver_array_0/in_13 subbyte2_wordline_driver_array_0/in_14 subbyte2_wordline_driver_array_0/in_15
+ subbyte2_wordline_driver_array_0/in_16 subbyte2_wordline_driver_array_0/in_17 subbyte2_wordline_driver_array_0/in_18
+ subbyte2_wordline_driver_array_0/in_19 subbyte2_wordline_driver_array_0/in_20 subbyte2_wordline_driver_array_0/in_21
+ subbyte2_wordline_driver_array_0/in_22 subbyte2_wordline_driver_array_0/in_23 subbyte2_wordline_driver_array_0/in_24
+ subbyte2_wordline_driver_array_0/in_25 subbyte2_wordline_driver_array_0/in_26 subbyte2_wordline_driver_array_0/in_27
+ subbyte2_wordline_driver_array_0/in_28 subbyte2_wordline_driver_array_0/in_29 subbyte2_wordline_driver_array_0/in_30
+ subbyte2_wordline_driver_array_0/in_31 subbyte2_wordline_driver_array_0/in_32 subbyte2_wordline_driver_array_0/in_33
+ subbyte2_wordline_driver_array_0/in_34 subbyte2_wordline_driver_array_0/in_35 subbyte2_wordline_driver_array_0/in_36
+ subbyte2_wordline_driver_array_0/in_37 subbyte2_wordline_driver_array_0/in_38 subbyte2_wordline_driver_array_0/in_39
+ subbyte2_wordline_driver_array_0/in_40 subbyte2_wordline_driver_array_0/in_41 subbyte2_wordline_driver_array_0/in_42
+ subbyte2_wordline_driver_array_0/in_43 subbyte2_wordline_driver_array_0/in_44 subbyte2_wordline_driver_array_0/in_45
+ subbyte2_wordline_driver_array_0/in_46 subbyte2_wordline_driver_array_0/in_47 subbyte2_wordline_driver_array_0/in_48
+ subbyte2_wordline_driver_array_0/in_49 subbyte2_wordline_driver_array_0/in_50 subbyte2_wordline_driver_array_0/in_51
+ subbyte2_wordline_driver_array_0/in_52 subbyte2_wordline_driver_array_0/in_53 subbyte2_wordline_driver_array_0/in_54
+ subbyte2_wordline_driver_array_0/in_55 subbyte2_wordline_driver_array_0/in_56 subbyte2_wordline_driver_array_0/in_57
+ subbyte2_wordline_driver_array_0/in_58 subbyte2_wordline_driver_array_0/in_59 subbyte2_wordline_driver_array_0/in_60
+ subbyte2_wordline_driver_array_0/in_61 subbyte2_wordline_driver_array_0/in_62 subbyte2_wordline_driver_array_0/in_63
+ vdd_uq7 vdd_uq6 vdd_uq8 vdd_uq9 vdd_uq13 vdd_uq11 vdd_uq17 vdd_uq16 vdd_uq18 vdd_uq1
+ vdd_uq3 gnd subbyte2_hierarchical_decoder
Xsubbyte2_wordline_driver_array_0 subbyte2_wordline_driver_array_0/in_0 subbyte2_wordline_driver_array_0/in_1
+ subbyte2_wordline_driver_array_0/in_2 subbyte2_wordline_driver_array_0/in_3 subbyte2_wordline_driver_array_0/in_4
+ subbyte2_wordline_driver_array_0/in_5 subbyte2_wordline_driver_array_0/in_6 subbyte2_wordline_driver_array_0/in_7
+ subbyte2_wordline_driver_array_0/in_8 subbyte2_wordline_driver_array_0/in_9 subbyte2_wordline_driver_array_0/in_10
+ subbyte2_wordline_driver_array_0/in_11 subbyte2_wordline_driver_array_0/in_12 subbyte2_wordline_driver_array_0/in_13
+ subbyte2_wordline_driver_array_0/in_14 subbyte2_wordline_driver_array_0/in_15 subbyte2_wordline_driver_array_0/in_16
+ subbyte2_wordline_driver_array_0/in_17 subbyte2_wordline_driver_array_0/in_18 subbyte2_wordline_driver_array_0/in_19
+ subbyte2_wordline_driver_array_0/in_20 subbyte2_wordline_driver_array_0/in_21 subbyte2_wordline_driver_array_0/in_22
+ subbyte2_wordline_driver_array_0/in_23 subbyte2_wordline_driver_array_0/in_24 subbyte2_wordline_driver_array_0/in_25
+ subbyte2_wordline_driver_array_0/in_26 subbyte2_wordline_driver_array_0/in_27 subbyte2_wordline_driver_array_0/in_28
+ subbyte2_wordline_driver_array_0/in_29 subbyte2_wordline_driver_array_0/in_30 subbyte2_wordline_driver_array_0/in_31
+ subbyte2_wordline_driver_array_0/in_32 subbyte2_wordline_driver_array_0/in_33 subbyte2_wordline_driver_array_0/in_34
+ subbyte2_wordline_driver_array_0/in_35 subbyte2_wordline_driver_array_0/in_36 subbyte2_wordline_driver_array_0/in_37
+ subbyte2_wordline_driver_array_0/in_38 subbyte2_wordline_driver_array_0/in_39 subbyte2_wordline_driver_array_0/in_40
+ subbyte2_wordline_driver_array_0/in_41 subbyte2_wordline_driver_array_0/in_42 subbyte2_wordline_driver_array_0/in_43
+ subbyte2_wordline_driver_array_0/in_44 subbyte2_wordline_driver_array_0/in_45 subbyte2_wordline_driver_array_0/in_46
+ subbyte2_wordline_driver_array_0/in_47 subbyte2_wordline_driver_array_0/in_48 subbyte2_wordline_driver_array_0/in_49
+ subbyte2_wordline_driver_array_0/in_50 subbyte2_wordline_driver_array_0/in_51 subbyte2_wordline_driver_array_0/in_52
+ subbyte2_wordline_driver_array_0/in_53 subbyte2_wordline_driver_array_0/in_54 subbyte2_wordline_driver_array_0/in_55
+ subbyte2_wordline_driver_array_0/in_56 subbyte2_wordline_driver_array_0/in_57 subbyte2_wordline_driver_array_0/in_58
+ subbyte2_wordline_driver_array_0/in_59 subbyte2_wordline_driver_array_0/in_60 subbyte2_wordline_driver_array_0/in_61
+ subbyte2_wordline_driver_array_0/in_62 subbyte2_wordline_driver_array_0/in_63 wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29
+ wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43
+ wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57
+ wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_en vdd vdd_uq0 gnd subbyte2_wordline_driver_array
.ends

.subckt subbyte2_pdriver A Z vdd gnd
Xsubbyte2_pinv_0 A Z vdd gnd subbyte2_pinv
.ends

.subckt subbyte2_pand2 A B Z gnd vdd
Xsubbyte2_pdriver_0 subbyte2_pnand2_0/Z Z vdd gnd subbyte2_pdriver
Xsubbyte2_pnand2_0 A B subbyte2_pnand2_0/Z vdd vdd gnd subbyte2_pnand2
.ends

.subckt subbyte2_hierarchical_predecode2x4_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd_uq0
+ gnd vdd
Xsubbyte2_pinv_0_0 in_1 subbyte2_pand2_3/B vdd_uq0 gnd subbyte2_pinv_0
Xsubbyte2_pinv_0_1 in_0 subbyte2_pand2_3/A vdd_uq0 gnd subbyte2_pinv_0
Xsubbyte2_pand2_0 in_0 in_1 out_3 gnd vdd subbyte2_pand2
Xsubbyte2_pand2_1 subbyte2_pand2_3/A in_1 out_2 gnd vdd subbyte2_pand2
Xsubbyte2_pand2_3 subbyte2_pand2_3/A subbyte2_pand2_3/B out_0 gnd vdd_uq0 subbyte2_pand2
Xsubbyte2_pand2_2 in_0 subbyte2_pand2_3/B out_1 gnd vdd_uq0 subbyte2_pand2
.ends

.subckt subbyte2_column_decoder in_0 in_1 out_0 out_1 out_2 out_3 gnd vdd
Xsubbyte2_hierarchical_predecode2x4_0_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
+ vdd subbyte2_hierarchical_predecode2x4_0
.ends

.subckt subbyte2_bank rbl_bl_0_0 rbl_bl_1_1 din0_6 din0_7 addr0_0 addr0_1 s_en1 p_en_bar0
+ w_en0 wl_en0 vdd_uq0 vdd_uq42 vdd_uq45 addr1_7 vdd_uq35 vdd_uq22 addr1_6 vdd_uq32
+ wl_en1 vdd_uq25 addr1_5 vdd_uq16 addr1_4 addr1_3 addr1_1 addr1_2 addr1_0 addr0_7
+ vdd_uq46 addr0_6 dout1_4 addr0_5 dout1_3 addr0_4 dout1_2 vdd_uq36 vdd_uq37 addr0_3
+ dout1_1 din0_5 vdd_uq43 addr0_2 dout1_0 vdd_uq26 vdd_uq44 din0_3 vdd_uq15 vdd_uq50
+ din0_2 vdd_uq17 din0_1 vdd_uq7 vdd_uq27 vdd_uq34 din0_4 vdd_uq12 dout1_7 din0_0
+ vdd_uq33 vdd_uq47 vdd_uq23 vdd_uq8 vdd_uq9 dout1_6 vdd_uq11 vdd_uq48 p_en_bar1 vdd_uq14
+ vdd_uq3 vdd_uq4 vdd_uq24 vdd_uq2 vdd dout1_5 vdd_uq6 vdd_uq49 vdd_uq13 gnd
Xsubbyte2_capped_replica_bitcell_array_0 rbl_bl_0_0 subbyte2_capped_replica_bitcell_array_0/rbl_bl_1_0
+ subbyte2_capped_replica_bitcell_array_0/rbl_br_1_0 subbyte2_port_data_0_0/br_0 subbyte2_port_data_0_0/br_1
+ subbyte2_port_data_0_0/br_2 subbyte2_port_data_0_0/br_3 subbyte2_port_data_0_0/bl_4
+ subbyte2_port_data_0_0/br_4 subbyte2_port_data_0_0/bl_5 subbyte2_port_data_0_0/br_5
+ subbyte2_port_data_0_0/bl_6 subbyte2_port_data_0_0/br_6 subbyte2_port_data_0_0/bl_7
+ subbyte2_port_data_0_0/br_7 subbyte2_port_data_0_0/bl_8 subbyte2_port_data_0_0/br_8
+ subbyte2_port_data_0_0/bl_9 subbyte2_port_data_0_0/bl_10 subbyte2_port_data_0_0/br_10
+ subbyte2_port_data_0_0/br_11 subbyte2_port_data_0_0/bl_12 subbyte2_port_data_0_0/br_12
+ subbyte2_port_data_0_0/bl_13 subbyte2_port_data_0_0/br_13 subbyte2_port_data_0_0/bl_14
+ subbyte2_port_data_0_0/br_14 subbyte2_port_data_0_0/bl_15 subbyte2_port_data_0_0/br_15
+ subbyte2_port_data_0_0/bl_16 subbyte2_port_data_0_0/br_16 subbyte2_port_data_0_0/bl_17
+ subbyte2_port_data_0_0/br_17 subbyte2_port_data_0_0/bl_18 subbyte2_port_data_0_0/br_18
+ subbyte2_port_data_0/bl_19 subbyte2_port_data_0_0/bl_19 subbyte2_port_data_0/br_19
+ subbyte2_port_data_0_0/bl_20 subbyte2_port_data_0_0/br_20 subbyte2_port_data_0_0/bl_21
+ subbyte2_port_data_0_0/br_21 subbyte2_port_data_0_0/br_22 subbyte2_port_data_0_0/bl_23
+ subbyte2_port_data_0_0/br_23 subbyte2_port_data_0_0/bl_24 subbyte2_port_data_0_0/br_24
+ subbyte2_port_data_0_0/bl_25 subbyte2_port_data_0_0/br_25 subbyte2_port_data_0_0/bl_26
+ subbyte2_port_data_0_0/br_26 subbyte2_port_data_0_0/bl_27 subbyte2_port_data_0_0/br_27
+ subbyte2_port_data_0_0/bl_28 subbyte2_port_data_0_0/br_28 subbyte2_port_data_0/bl_29
+ subbyte2_port_data_0_0/bl_29 subbyte2_port_data_0/bl_30 subbyte2_port_data_0_0/bl_30
+ subbyte2_port_data_0_0/br_30 subbyte2_port_data_0_0/bl_31 subbyte2_port_data_0_0/br_31
+ subbyte2_capped_replica_bitcell_array_0/rbl_bl_0_1 rbl_bl_1_1 subbyte2_capped_replica_bitcell_array_0/rbl_br_0_1
+ subbyte2_port_address_0/rbl_wl subbyte2_port_address_0/wl_1 subbyte2_port_address_0/wl_2
+ subbyte2_port_address_0/wl_3 subbyte2_port_address_0/wl_4 subbyte2_port_address_0/wl_5
+ subbyte2_port_address_0/wl_6 subbyte2_port_address_0/wl_7 subbyte2_port_address_0/wl_8
+ subbyte2_port_address_0_0/wl_10 subbyte2_port_address_0_0/wl_11 subbyte2_port_address_0_0/wl_12
+ subbyte2_port_address_0_0/wl_13 subbyte2_port_address_0_0/wl_14 subbyte2_port_address_0/wl_15
+ subbyte2_port_address_0_0/wl_15 subbyte2_port_address_0/wl_16 subbyte2_port_address_0_0/wl_16
+ subbyte2_port_address_0/wl_17 subbyte2_port_address_0_0/wl_17 subbyte2_port_address_0/wl_18
+ subbyte2_port_address_0_0/wl_18 subbyte2_port_address_0_0/wl_19 subbyte2_port_address_0_0/wl_20
+ subbyte2_port_address_0_0/wl_21 subbyte2_port_address_0_0/wl_22 subbyte2_port_address_0_0/wl_23
+ subbyte2_port_address_0_0/wl_24 subbyte2_port_address_0_0/wl_25 subbyte2_port_address_0/wl_26
+ subbyte2_port_address_0_0/wl_26 subbyte2_port_address_0/wl_27 subbyte2_port_address_0_0/wl_27
+ subbyte2_port_address_0/wl_28 subbyte2_port_address_0_0/wl_28 subbyte2_port_address_0_0/wl_29
+ subbyte2_port_address_0_0/wl_30 subbyte2_port_address_0_0/wl_31 subbyte2_port_address_0_0/wl_32
+ subbyte2_port_address_0_0/wl_33 subbyte2_port_address_0_0/wl_34 subbyte2_port_address_0_0/wl_35
+ subbyte2_port_address_0_0/wl_36 subbyte2_port_address_0/wl_37 subbyte2_port_address_0_0/wl_37
+ subbyte2_port_address_0/wl_38 subbyte2_port_address_0_0/wl_38 subbyte2_port_address_0_0/wl_39
+ subbyte2_port_address_0_0/wl_40 subbyte2_port_address_0_0/wl_41 subbyte2_port_address_0_0/wl_42
+ subbyte2_port_address_0_0/wl_43 subbyte2_port_address_0_0/wl_44 subbyte2_port_address_0_0/wl_45
+ subbyte2_port_address_0_0/wl_46 subbyte2_port_address_0_0/wl_47 subbyte2_port_address_0/wl_48
+ subbyte2_port_address_0_0/wl_48 subbyte2_port_address_0/wl_49 subbyte2_port_address_0_0/wl_49
+ subbyte2_port_address_0_0/wl_50 subbyte2_port_address_0_0/wl_51 subbyte2_port_address_0_0/wl_52
+ subbyte2_port_address_0_0/wl_53 subbyte2_port_address_0_0/wl_54 subbyte2_port_address_0_0/wl_55
+ subbyte2_port_address_0_0/wl_56 subbyte2_port_address_0_0/wl_57 subbyte2_port_address_0_0/wl_58
+ subbyte2_port_address_0/wl_59 subbyte2_port_address_0_0/wl_59 subbyte2_port_address_0/wl_60
+ subbyte2_port_address_0_0/wl_60 subbyte2_port_address_0_0/wl_61 subbyte2_port_address_0_0/wl_62
+ subbyte2_port_address_0_0/wl_63 subbyte2_port_address_0_0/rbl_wl subbyte2_port_address_0_0/wl_9
+ subbyte2_port_address_0_0/wl_8 subbyte2_port_address_0_0/wl_7 subbyte2_port_address_0_0/wl_6
+ subbyte2_port_data_0/br_8 subbyte2_port_address_0_0/wl_5 subbyte2_port_data_0/br_7
+ subbyte2_port_data_0/br_18 subbyte2_port_data_0/bl_8 subbyte2_port_address_0_0/wl_4
+ subbyte2_port_data_0/br_6 subbyte2_port_data_0/br_17 subbyte2_port_data_0/br_28
+ subbyte2_port_data_0/bl_7 subbyte2_port_address_0_0/wl_3 subbyte2_port_data_0/br_5
+ subbyte2_port_data_0/br_16 subbyte2_port_data_0/br_27 subbyte2_port_data_0/bl_6
+ subbyte2_port_address_0_0/wl_2 subbyte2_port_data_0/br_4 subbyte2_port_data_0/br_15
+ subbyte2_port_data_0/br_26 subbyte2_port_data_0/bl_5 subbyte2_port_address_0_0/wl_1
+ subbyte2_port_data_0/br_3 subbyte2_port_data_0/br_25 subbyte2_port_data_0/br_14
+ subbyte2_port_data_0/bl_4 subbyte2_port_address_0_0/wl_0 subbyte2_port_data_0/br_2
+ subbyte2_port_data_0/br_13 subbyte2_port_data_0/br_24 subbyte2_port_data_0/bl_3
+ subbyte2_port_data_0/br_1 subbyte2_port_data_0/bl_18 subbyte2_port_data_0/br_23
+ subbyte2_port_data_0/br_12 subbyte2_port_data_0/bl_2 subbyte2_port_data_0/bl_17
+ subbyte2_port_data_0/bl_28 subbyte2_port_address_0/wl_25 subbyte2_port_address_0/wl_14
+ subbyte2_port_data_0/br_0 subbyte2_port_address_0/wl_58 subbyte2_port_address_0/wl_47
+ subbyte2_port_address_0/wl_36 subbyte2_port_data_0/br_11 subbyte2_port_data_0/br_22
+ subbyte2_port_data_0/bl_1 subbyte2_port_data_0/bl_16 subbyte2_port_data_0/bl_27
+ subbyte2_port_address_0/wl_46 subbyte2_port_address_0/wl_35 subbyte2_port_address_0/wl_13
+ subbyte2_port_address_0/wl_24 subbyte2_port_data_0/rbl_br subbyte2_port_address_0/wl_57
+ subbyte2_port_data_0/br_10 subbyte2_port_data_0/br_21 subbyte2_port_data_0/bl_0
+ subbyte2_port_data_0_0/bl_3 subbyte2_port_data_0/bl_26 subbyte2_port_address_0/wl_34
+ subbyte2_port_address_0/wl_23 subbyte2_port_address_0/wl_56 subbyte2_port_address_0/wl_12
+ subbyte2_port_address_0/wl_45 subbyte2_port_data_0/bl_15 subbyte2_port_data_0/br_31
+ subbyte2_port_data_0/br_20 subbyte2_port_data_0/br_9 subbyte2_port_data_0_0/bl_2
+ subbyte2_port_data_0/bl_25 subbyte2_port_data_0/bl_14 subbyte2_port_address_0/wl_11
+ subbyte2_port_address_0/wl_55 subbyte2_port_address_0/wl_22 subbyte2_port_address_0/wl_33
+ subbyte2_port_address_0/wl_44 subbyte2_port_data_0/br_30 subbyte2_port_data_0_0/rbl_br
+ subbyte2_port_data_0_0/bl_1 subbyte2_port_data_0/bl_24 subbyte2_port_data_0/bl_13
+ subbyte2_port_address_0/wl_54 subbyte2_port_address_0/wl_43 subbyte2_port_address_0/wl_32
+ subbyte2_port_address_0/wl_21 subbyte2_port_address_0/wl_10 subbyte2_port_data_0/br_29
+ subbyte2_port_data_0_0/br_9 subbyte2_port_data_0_0/bl_0 subbyte2_port_address_0/wl_0
+ subbyte2_port_data_0/bl_12 subbyte2_port_data_0/bl_23 subbyte2_port_address_0/wl_31
+ subbyte2_port_address_0/wl_42 subbyte2_port_address_0/wl_9 subbyte2_port_address_0/wl_20
+ subbyte2_port_address_0/wl_53 subbyte2_port_data_0_0/br_19 subbyte2_port_data_0/bl_11
+ subbyte2_port_data_0/bl_22 subbyte2_port_address_0/wl_63 subbyte2_port_address_0/wl_30
+ subbyte2_port_address_0/wl_19 subbyte2_port_address_0/wl_41 subbyte2_port_address_0/wl_52
+ subbyte2_port_data_0_0/br_29 subbyte2_port_address_0/wl_62 subbyte2_port_address_0/wl_51
+ subbyte2_port_data_0/bl_10 subbyte2_port_data_0/bl_21 subbyte2_port_address_0/wl_29
+ subbyte2_port_address_0/wl_40 subbyte2_port_data_0/bl_9 subbyte2_port_address_0/wl_50
+ subbyte2_port_address_0/wl_39 subbyte2_port_data_0/bl_31 subbyte2_port_data_0/bl_20
+ subbyte2_port_address_0/wl_61 subbyte2_port_data_0_0/bl_11 subbyte2_port_data_0_0/bl_22
+ vdd_uq6 gnd subbyte2_capped_replica_bitcell_array
Xsubbyte2_port_data_0_0 rbl_bl_1_1 subbyte2_port_data_0_0/rbl_br subbyte2_port_data_0_0/bl_0
+ subbyte2_port_data_0_0/br_0 subbyte2_port_data_0_0/bl_1 subbyte2_port_data_0_0/br_1
+ subbyte2_port_data_0_0/bl_2 subbyte2_port_data_0_0/br_2 subbyte2_port_data_0_0/bl_3
+ subbyte2_port_data_0_0/br_3 subbyte2_port_data_0_0/bl_4 subbyte2_port_data_0_0/br_4
+ subbyte2_port_data_0_0/bl_5 subbyte2_port_data_0_0/br_5 subbyte2_port_data_0_0/bl_6
+ subbyte2_port_data_0_0/br_6 subbyte2_port_data_0_0/bl_7 subbyte2_port_data_0_0/br_7
+ subbyte2_port_data_0_0/bl_8 subbyte2_port_data_0_0/br_8 subbyte2_port_data_0_0/bl_9
+ subbyte2_port_data_0_0/br_9 subbyte2_port_data_0_0/bl_10 subbyte2_port_data_0_0/br_10
+ subbyte2_port_data_0_0/bl_11 subbyte2_port_data_0_0/br_11 subbyte2_port_data_0_0/bl_12
+ subbyte2_port_data_0_0/br_12 subbyte2_port_data_0_0/bl_13 subbyte2_port_data_0_0/br_13
+ subbyte2_port_data_0_0/bl_14 subbyte2_port_data_0_0/br_14 subbyte2_port_data_0_0/bl_15
+ subbyte2_port_data_0_0/br_15 subbyte2_port_data_0_0/bl_16 subbyte2_port_data_0_0/br_16
+ subbyte2_port_data_0_0/bl_17 subbyte2_port_data_0_0/br_17 subbyte2_port_data_0_0/bl_18
+ subbyte2_port_data_0_0/br_18 subbyte2_port_data_0_0/bl_19 subbyte2_port_data_0_0/br_19
+ subbyte2_port_data_0_0/bl_20 subbyte2_port_data_0_0/br_20 subbyte2_port_data_0_0/bl_21
+ subbyte2_port_data_0_0/br_21 subbyte2_port_data_0_0/bl_22 subbyte2_port_data_0_0/br_22
+ subbyte2_port_data_0_0/bl_23 subbyte2_port_data_0_0/br_23 subbyte2_port_data_0_0/bl_24
+ subbyte2_port_data_0_0/br_24 subbyte2_port_data_0_0/bl_25 subbyte2_port_data_0_0/br_25
+ subbyte2_port_data_0_0/bl_26 subbyte2_port_data_0_0/br_26 subbyte2_port_data_0_0/bl_27
+ subbyte2_port_data_0_0/br_27 subbyte2_port_data_0_0/bl_28 subbyte2_port_data_0_0/br_28
+ subbyte2_port_data_0_0/bl_29 subbyte2_port_data_0_0/br_29 subbyte2_port_data_0_0/bl_30
+ subbyte2_port_data_0_0/br_30 subbyte2_port_data_0_0/bl_31 subbyte2_port_data_0_0/br_31
+ dout1_1 dout1_2 dout1_5 dout1_6 subbyte2_port_data_0_0/sel_3 vdd_uq48 dout1_4 subbyte2_port_data_0_0/sel_2
+ subbyte2_port_data_0_0/sel_1 s_en1 dout1_0 subbyte2_port_data_0_0/sel_0 dout1_3
+ vdd_uq50 vdd_uq49 dout1_7 p_en_bar1 gnd subbyte2_port_data_0
Xsubbyte2_port_data_0 rbl_bl_0_0 subbyte2_port_data_0/rbl_br subbyte2_port_data_0/bl_0
+ subbyte2_port_data_0/br_0 subbyte2_port_data_0/bl_1 subbyte2_port_data_0/br_1 subbyte2_port_data_0/bl_2
+ subbyte2_port_data_0/br_2 subbyte2_port_data_0/bl_3 subbyte2_port_data_0/br_3 subbyte2_port_data_0/bl_4
+ subbyte2_port_data_0/br_4 subbyte2_port_data_0/bl_5 subbyte2_port_data_0/br_5 subbyte2_port_data_0/bl_6
+ subbyte2_port_data_0/br_6 subbyte2_port_data_0/bl_7 subbyte2_port_data_0/br_7 subbyte2_port_data_0/bl_8
+ subbyte2_port_data_0/br_8 subbyte2_port_data_0/bl_9 subbyte2_port_data_0/br_9 subbyte2_port_data_0/bl_10
+ subbyte2_port_data_0/br_10 subbyte2_port_data_0/bl_11 subbyte2_port_data_0/br_11
+ subbyte2_port_data_0/bl_12 subbyte2_port_data_0/br_12 subbyte2_port_data_0/bl_13
+ subbyte2_port_data_0/br_13 subbyte2_port_data_0/bl_14 subbyte2_port_data_0/br_14
+ subbyte2_port_data_0/bl_15 subbyte2_port_data_0/br_15 subbyte2_port_data_0/bl_16
+ subbyte2_port_data_0/br_16 subbyte2_port_data_0/bl_17 subbyte2_port_data_0/br_17
+ subbyte2_port_data_0/bl_18 subbyte2_port_data_0/br_18 subbyte2_port_data_0/bl_19
+ subbyte2_port_data_0/br_19 subbyte2_port_data_0/bl_20 subbyte2_port_data_0/br_20
+ subbyte2_port_data_0/bl_21 subbyte2_port_data_0/br_21 subbyte2_port_data_0/bl_22
+ subbyte2_port_data_0/br_22 subbyte2_port_data_0/bl_23 subbyte2_port_data_0/br_23
+ subbyte2_port_data_0/bl_24 subbyte2_port_data_0/br_24 subbyte2_port_data_0/bl_25
+ subbyte2_port_data_0/br_25 subbyte2_port_data_0/bl_26 subbyte2_port_data_0/br_26
+ subbyte2_port_data_0/bl_27 subbyte2_port_data_0/br_27 subbyte2_port_data_0/bl_28
+ subbyte2_port_data_0/br_28 subbyte2_port_data_0/bl_29 subbyte2_port_data_0/br_29
+ subbyte2_port_data_0/bl_30 subbyte2_port_data_0/br_30 subbyte2_port_data_0/bl_31
+ subbyte2_port_data_0/br_31 din0_7 subbyte2_port_data_0/sel_3 din0_2 din0_1 din0_4
+ din0_5 subbyte2_port_data_0/sel_2 subbyte2_port_data_0/sel_1 subbyte2_port_data_0/sel_0
+ w_en0 din0_0 din0_3 p_en_bar0 vdd_uq14 din0_6 vdd_uq13 vdd_uq15 gnd subbyte2_port_data
Xsubbyte2_port_address_0 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 wl_en0 subbyte2_port_address_0/wl_0
+ subbyte2_port_address_0/wl_1 subbyte2_port_address_0/wl_2 subbyte2_port_address_0/wl_3
+ subbyte2_port_address_0/wl_4 subbyte2_port_address_0/wl_5 subbyte2_port_address_0/wl_6
+ subbyte2_port_address_0/wl_7 subbyte2_port_address_0/wl_8 subbyte2_port_address_0/wl_9
+ subbyte2_port_address_0/wl_10 subbyte2_port_address_0/wl_11 subbyte2_port_address_0/wl_12
+ subbyte2_port_address_0/wl_13 subbyte2_port_address_0/wl_14 subbyte2_port_address_0/wl_15
+ subbyte2_port_address_0/wl_16 subbyte2_port_address_0/wl_17 subbyte2_port_address_0/wl_18
+ subbyte2_port_address_0/wl_19 subbyte2_port_address_0/wl_20 subbyte2_port_address_0/wl_21
+ subbyte2_port_address_0/wl_22 subbyte2_port_address_0/wl_23 subbyte2_port_address_0/wl_24
+ subbyte2_port_address_0/wl_25 subbyte2_port_address_0/wl_26 subbyte2_port_address_0/wl_27
+ subbyte2_port_address_0/wl_28 subbyte2_port_address_0/wl_29 subbyte2_port_address_0/wl_30
+ subbyte2_port_address_0/wl_31 subbyte2_port_address_0/wl_32 subbyte2_port_address_0/wl_33
+ subbyte2_port_address_0/wl_34 subbyte2_port_address_0/wl_35 subbyte2_port_address_0/wl_36
+ subbyte2_port_address_0/wl_37 subbyte2_port_address_0/wl_38 subbyte2_port_address_0/wl_39
+ subbyte2_port_address_0/wl_40 subbyte2_port_address_0/wl_41 subbyte2_port_address_0/wl_42
+ subbyte2_port_address_0/wl_43 subbyte2_port_address_0/wl_44 subbyte2_port_address_0/wl_45
+ subbyte2_port_address_0/wl_46 subbyte2_port_address_0/wl_47 subbyte2_port_address_0/wl_48
+ subbyte2_port_address_0/wl_49 subbyte2_port_address_0/wl_50 subbyte2_port_address_0/wl_51
+ subbyte2_port_address_0/wl_52 subbyte2_port_address_0/wl_53 subbyte2_port_address_0/wl_54
+ subbyte2_port_address_0/wl_55 subbyte2_port_address_0/wl_56 subbyte2_port_address_0/wl_57
+ subbyte2_port_address_0/wl_58 subbyte2_port_address_0/wl_59 subbyte2_port_address_0/wl_60
+ subbyte2_port_address_0/wl_61 subbyte2_port_address_0/wl_62 subbyte2_port_address_0/wl_63
+ subbyte2_port_address_0/rbl_wl vdd_uq25 vdd_uq26 vdd_uq22 vdd_uq16 vdd_uq45 vdd_uq42
+ vdd_uq32 vdd_uq35 vdd_uq36 vdd_uq46 vdd_uq7 vdd_uq8 vdd_uq11 vdd_uq9 gnd subbyte2_port_address
Xsubbyte2_port_address_0_0 addr1_2 addr1_3 addr1_4 addr1_5 addr1_6 addr1_7 wl_en1
+ subbyte2_port_address_0_0/wl_0 subbyte2_port_address_0_0/wl_1 subbyte2_port_address_0_0/wl_2
+ subbyte2_port_address_0_0/wl_3 subbyte2_port_address_0_0/wl_4 subbyte2_port_address_0_0/wl_5
+ subbyte2_port_address_0_0/wl_6 subbyte2_port_address_0_0/wl_7 subbyte2_port_address_0_0/wl_8
+ subbyte2_port_address_0_0/wl_9 subbyte2_port_address_0_0/wl_10 subbyte2_port_address_0_0/wl_11
+ subbyte2_port_address_0_0/wl_12 subbyte2_port_address_0_0/wl_13 subbyte2_port_address_0_0/wl_14
+ subbyte2_port_address_0_0/wl_15 subbyte2_port_address_0_0/wl_16 subbyte2_port_address_0_0/wl_17
+ subbyte2_port_address_0_0/wl_18 subbyte2_port_address_0_0/wl_19 subbyte2_port_address_0_0/wl_20
+ subbyte2_port_address_0_0/wl_21 subbyte2_port_address_0_0/wl_22 subbyte2_port_address_0_0/wl_23
+ subbyte2_port_address_0_0/wl_24 subbyte2_port_address_0_0/wl_25 subbyte2_port_address_0_0/wl_26
+ subbyte2_port_address_0_0/wl_27 subbyte2_port_address_0_0/wl_28 subbyte2_port_address_0_0/wl_29
+ subbyte2_port_address_0_0/wl_30 subbyte2_port_address_0_0/wl_31 subbyte2_port_address_0_0/wl_32
+ subbyte2_port_address_0_0/wl_33 subbyte2_port_address_0_0/wl_34 subbyte2_port_address_0_0/wl_35
+ subbyte2_port_address_0_0/wl_36 subbyte2_port_address_0_0/wl_37 subbyte2_port_address_0_0/wl_38
+ subbyte2_port_address_0_0/wl_39 subbyte2_port_address_0_0/wl_40 subbyte2_port_address_0_0/wl_41
+ subbyte2_port_address_0_0/wl_42 subbyte2_port_address_0_0/wl_43 subbyte2_port_address_0_0/wl_44
+ subbyte2_port_address_0_0/wl_45 subbyte2_port_address_0_0/wl_46 subbyte2_port_address_0_0/wl_47
+ subbyte2_port_address_0_0/wl_48 subbyte2_port_address_0_0/wl_49 subbyte2_port_address_0_0/wl_50
+ subbyte2_port_address_0_0/wl_51 subbyte2_port_address_0_0/wl_52 subbyte2_port_address_0_0/wl_53
+ subbyte2_port_address_0_0/wl_54 subbyte2_port_address_0_0/wl_55 subbyte2_port_address_0_0/wl_56
+ subbyte2_port_address_0_0/wl_57 subbyte2_port_address_0_0/wl_58 subbyte2_port_address_0_0/wl_59
+ subbyte2_port_address_0_0/wl_60 subbyte2_port_address_0_0/wl_61 subbyte2_port_address_0_0/wl_62
+ subbyte2_port_address_0_0/wl_63 subbyte2_port_address_0_0/rbl_wl vdd vdd_uq24 vdd_uq23
+ vdd_uq17 vdd_uq47 vdd_uq44 vdd_uq37 vdd_uq27 vdd_uq34 vdd_uq33 vdd_uq43 vdd_uq4
+ vdd_uq3 gnd vdd_uq2 subbyte2_port_address_0
Xsubbyte2_column_decoder_0 addr1_0 addr1_1 subbyte2_port_data_0_0/sel_0 subbyte2_port_data_0_0/sel_1
+ subbyte2_port_data_0_0/sel_2 subbyte2_port_data_0_0/sel_3 gnd vdd_uq12 subbyte2_column_decoder
Xsubbyte2_column_decoder_1 addr0_0 addr0_1 subbyte2_port_data_0/sel_0 subbyte2_port_data_0/sel_1
+ subbyte2_port_data_0/sel_2 subbyte2_port_data_0/sel_3 gnd vdd_uq0 subbyte2_column_decoder
.ends

.subckt subbyte2_col_addr_dff dout_0 dout_1 clk din_0 vdd gnd din_1
Xsky130_fd_bd_sram__openram_dff_0 din_1 dout_1 gnd clk vdd sky130_fd_bd_sram__openram_dff_0/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 din_0 dout_0 gnd clk vdd sky130_fd_bd_sram__openram_dff_1/QN
+ sky130_fd_bd_sram__openram_dff
.ends

.subckt subbyte2_row_addr_dff din_1 dout_0 dout_2 dout_4 clk din_4 dout_5 din_2 din_0
+ dout_3 dout_1 gnd din_5 din_3 vdd
Xsky130_fd_bd_sram__openram_dff_5 din_0 dout_0 gnd clk vdd sky130_fd_bd_sram__openram_dff_5/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_0 din_5 dout_5 gnd clk vdd sky130_fd_bd_sram__openram_dff_0/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 din_4 dout_4 gnd clk vdd sky130_fd_bd_sram__openram_dff_1/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_2 din_3 dout_3 gnd clk vdd sky130_fd_bd_sram__openram_dff_2/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_4 din_1 dout_1 gnd clk vdd sky130_fd_bd_sram__openram_dff_4/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_3 din_2 dout_2 gnd clk vdd sky130_fd_bd_sram__openram_dff_3/QN
+ sky130_fd_bd_sram__openram_dff
.ends

.subckt subbyte2_data_dff din_1 din_3 din_7 dout_0 dout_2 dout_4 dout_6 clk vdd din_6
+ din_4 dout_7 dout_5 din_2 din_0 dout_3 dout_1 gnd din_5
Xsky130_fd_bd_sram__openram_dff_5 din_2 dout_2 gnd clk vdd sky130_fd_bd_sram__openram_dff_5/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_6 din_1 dout_1 gnd clk vdd sky130_fd_bd_sram__openram_dff_6/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_7 din_0 dout_0 gnd clk vdd sky130_fd_bd_sram__openram_dff_7/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_0 din_7 dout_7 gnd clk vdd sky130_fd_bd_sram__openram_dff_0/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_1 din_6 dout_6 gnd clk vdd sky130_fd_bd_sram__openram_dff_1/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_2 din_5 dout_5 gnd clk vdd sky130_fd_bd_sram__openram_dff_2/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_4 din_3 dout_3 gnd clk vdd sky130_fd_bd_sram__openram_dff_4/QN
+ sky130_fd_bd_sram__openram_dff
Xsky130_fd_bd_sram__openram_dff_3 din_4 dout_4 gnd clk vdd sky130_fd_bd_sram__openram_dff_3/QN
+ sky130_fd_bd_sram__openram_dff
.ends

.subckt subbyte2 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1]
+ addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 clk0 clk1 dout1[0]
+ dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] vccd1 vssd1
Xsubbyte2_control_logic_r_0 clk1 subbyte2_bank_0/rbl_bl_1_1 subbyte2_bank_0/s_en1
+ subbyte2_bank_0/p_en_bar1 subbyte2_bank_0/wl_en1 subbyte2_row_addr_dff_0/clk vccd1
+ csb1 vccd1 vssd1 vccd1 subbyte2_control_logic_r
Xsubbyte2_control_logic_w_0 clk0 subbyte2_bank_0/rbl_bl_0_0 subbyte2_bank_0/w_en0
+ subbyte2_bank_0/p_en_bar0 subbyte2_bank_0/wl_en0 subbyte2_data_dff_0/clk vccd1 csb0
+ vssd1 vccd1 vccd1 subbyte2_control_logic_w
Xsubbyte2_bank_0 subbyte2_bank_0/rbl_bl_0_0 subbyte2_bank_0/rbl_bl_1_1 subbyte2_bank_0/din0_6
+ subbyte2_bank_0/din0_7 subbyte2_bank_0/addr0_0 subbyte2_bank_0/addr0_1 subbyte2_bank_0/s_en1
+ subbyte2_bank_0/p_en_bar0 subbyte2_bank_0/w_en0 subbyte2_bank_0/wl_en0 vccd1 vccd1
+ vccd1 subbyte2_bank_0/addr1_7 vccd1 vccd1 subbyte2_bank_0/addr1_6 vccd1 subbyte2_bank_0/wl_en1
+ vccd1 subbyte2_bank_0/addr1_5 vccd1 subbyte2_bank_0/addr1_4 subbyte2_bank_0/addr1_3
+ subbyte2_bank_0/addr1_1 subbyte2_bank_0/addr1_2 subbyte2_bank_0/addr1_0 subbyte2_bank_0/addr0_7
+ vccd1 subbyte2_bank_0/addr0_6 dout1[4] subbyte2_bank_0/addr0_5 dout1[3] subbyte2_bank_0/addr0_4
+ dout1[2] vccd1 vccd1 subbyte2_bank_0/addr0_3 dout1[1] subbyte2_bank_0/din0_5 vccd1
+ subbyte2_bank_0/addr0_2 dout1[0] vccd1 vccd1 subbyte2_bank_0/din0_3 vccd1 vccd1
+ subbyte2_bank_0/din0_2 vccd1 subbyte2_bank_0/din0_1 vccd1 vccd1 vccd1 subbyte2_bank_0/din0_4
+ vccd1 dout1[7] subbyte2_bank_0/din0_0 vccd1 vccd1 vccd1 vccd1 vccd1 dout1[6] vccd1
+ vccd1 subbyte2_bank_0/p_en_bar1 vccd1 vccd1 vccd1 vccd1 vccd1 vccd1 dout1[5] vccd1
+ vccd1 vccd1 vssd1 subbyte2_bank
Xsubbyte2_col_addr_dff_0 subbyte2_bank_0/addr1_0 subbyte2_bank_0/addr1_1 subbyte2_row_addr_dff_0/clk
+ addr1[0] vccd1 vssd1 addr1[1] subbyte2_col_addr_dff
Xsubbyte2_col_addr_dff_1 subbyte2_bank_0/addr0_0 subbyte2_bank_0/addr0_1 subbyte2_data_dff_0/clk
+ addr0[0] vccd1 vssd1 addr0[1] subbyte2_col_addr_dff
Xsubbyte2_row_addr_dff_0 addr1[3] subbyte2_bank_0/addr1_2 subbyte2_bank_0/addr1_4
+ subbyte2_bank_0/addr1_6 subbyte2_row_addr_dff_0/clk addr1[6] subbyte2_bank_0/addr1_7
+ addr1[4] addr1[2] subbyte2_bank_0/addr1_5 subbyte2_bank_0/addr1_3 vssd1 addr1[7]
+ addr1[5] vccd1 subbyte2_row_addr_dff
Xsubbyte2_row_addr_dff_1 addr0[3] subbyte2_bank_0/addr0_2 subbyte2_bank_0/addr0_4
+ subbyte2_bank_0/addr0_6 subbyte2_data_dff_0/clk addr0[6] subbyte2_bank_0/addr0_7
+ addr0[4] addr0[2] subbyte2_bank_0/addr0_5 subbyte2_bank_0/addr0_3 vssd1 addr0[7]
+ addr0[5] vccd1 subbyte2_row_addr_dff
Xsubbyte2_data_dff_0 din0[1] din0[3] din0[7] subbyte2_bank_0/din0_0 subbyte2_bank_0/din0_2
+ subbyte2_bank_0/din0_4 subbyte2_bank_0/din0_6 subbyte2_data_dff_0/clk vccd1 din0[6]
+ din0[4] subbyte2_bank_0/din0_7 subbyte2_bank_0/din0_5 din0[2] din0[0] subbyte2_bank_0/din0_3
+ subbyte2_bank_0/din0_1 vssd1 din0[5] subbyte2_data_dff
.ends

