magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1260 -1173 23147 3444
<< poly >>
rect 2216 435 2246 896
rect 2840 559 2870 896
rect 3464 683 3494 896
rect 4088 807 4118 896
rect 4056 791 4122 807
rect 4056 757 4072 791
rect 4106 757 4122 791
rect 4056 741 4122 757
rect 3460 667 3526 683
rect 3460 633 3476 667
rect 3510 633 3526 667
rect 3460 617 3526 633
rect 2808 543 2874 559
rect 2808 509 2824 543
rect 2858 509 2874 543
rect 2808 493 2874 509
rect 4712 435 4742 896
rect 5336 559 5366 896
rect 5960 683 5990 896
rect 6584 807 6614 896
rect 6552 791 6618 807
rect 6552 757 6568 791
rect 6602 757 6618 791
rect 6552 741 6618 757
rect 5956 667 6022 683
rect 5956 633 5972 667
rect 6006 633 6022 667
rect 5956 617 6022 633
rect 5304 543 5370 559
rect 5304 509 5320 543
rect 5354 509 5370 543
rect 5304 493 5370 509
rect 7208 435 7238 896
rect 7832 559 7862 896
rect 8456 683 8486 896
rect 9080 807 9110 896
rect 9048 791 9114 807
rect 9048 757 9064 791
rect 9098 757 9114 791
rect 9048 741 9114 757
rect 8452 667 8518 683
rect 8452 633 8468 667
rect 8502 633 8518 667
rect 8452 617 8518 633
rect 7800 543 7866 559
rect 7800 509 7816 543
rect 7850 509 7866 543
rect 7800 493 7866 509
rect 9704 435 9734 896
rect 10328 559 10358 896
rect 10952 683 10982 896
rect 11576 807 11606 896
rect 11544 791 11610 807
rect 11544 757 11560 791
rect 11594 757 11610 791
rect 11544 741 11610 757
rect 10948 667 11014 683
rect 10948 633 10964 667
rect 10998 633 11014 667
rect 10948 617 11014 633
rect 10296 543 10362 559
rect 10296 509 10312 543
rect 10346 509 10362 543
rect 10296 493 10362 509
rect 12200 435 12230 896
rect 12824 559 12854 896
rect 13448 683 13478 896
rect 14072 807 14102 896
rect 14040 791 14106 807
rect 14040 757 14056 791
rect 14090 757 14106 791
rect 14040 741 14106 757
rect 13444 667 13510 683
rect 13444 633 13460 667
rect 13494 633 13510 667
rect 13444 617 13510 633
rect 12792 543 12858 559
rect 12792 509 12808 543
rect 12842 509 12858 543
rect 12792 493 12858 509
rect 14696 435 14726 896
rect 15320 559 15350 896
rect 15944 683 15974 896
rect 16568 807 16598 896
rect 16536 791 16602 807
rect 16536 757 16552 791
rect 16586 757 16602 791
rect 16536 741 16602 757
rect 15940 667 16006 683
rect 15940 633 15956 667
rect 15990 633 16006 667
rect 15940 617 16006 633
rect 15288 543 15354 559
rect 15288 509 15304 543
rect 15338 509 15354 543
rect 15288 493 15354 509
rect 17192 435 17222 896
rect 17816 559 17846 896
rect 18440 683 18470 896
rect 19064 807 19094 896
rect 19032 791 19098 807
rect 19032 757 19048 791
rect 19082 757 19098 791
rect 19032 741 19098 757
rect 18436 667 18502 683
rect 18436 633 18452 667
rect 18486 633 18502 667
rect 18436 617 18502 633
rect 17784 543 17850 559
rect 17784 509 17800 543
rect 17834 509 17850 543
rect 17784 493 17850 509
rect 19688 435 19718 896
rect 20312 559 20342 896
rect 20936 683 20966 896
rect 21560 807 21590 896
rect 21528 791 21594 807
rect 21528 757 21544 791
rect 21578 757 21594 791
rect 21528 741 21594 757
rect 20932 667 20998 683
rect 20932 633 20948 667
rect 20982 633 20998 667
rect 20932 617 20998 633
rect 20280 543 20346 559
rect 20280 509 20296 543
rect 20330 509 20346 543
rect 20280 493 20346 509
rect 2212 419 2278 435
rect 2212 385 2228 419
rect 2262 385 2278 419
rect 2212 369 2278 385
rect 4708 419 4774 435
rect 4708 385 4724 419
rect 4758 385 4774 419
rect 4708 369 4774 385
rect 7204 419 7270 435
rect 7204 385 7220 419
rect 7254 385 7270 419
rect 7204 369 7270 385
rect 9700 419 9766 435
rect 9700 385 9716 419
rect 9750 385 9766 419
rect 9700 369 9766 385
rect 12196 419 12262 435
rect 12196 385 12212 419
rect 12246 385 12262 419
rect 12196 369 12262 385
rect 14692 419 14758 435
rect 14692 385 14708 419
rect 14742 385 14758 419
rect 14692 369 14758 385
rect 17188 419 17254 435
rect 17188 385 17204 419
rect 17238 385 17254 419
rect 17188 369 17254 385
rect 19684 419 19750 435
rect 19684 385 19700 419
rect 19734 385 19750 419
rect 19684 369 19750 385
<< polycont >>
rect 4072 757 4106 791
rect 3476 633 3510 667
rect 2824 509 2858 543
rect 6568 757 6602 791
rect 5972 633 6006 667
rect 5320 509 5354 543
rect 9064 757 9098 791
rect 8468 633 8502 667
rect 7816 509 7850 543
rect 11560 757 11594 791
rect 10964 633 10998 667
rect 10312 509 10346 543
rect 14056 757 14090 791
rect 13460 633 13494 667
rect 12808 509 12842 543
rect 16552 757 16586 791
rect 15956 633 15990 667
rect 15304 509 15338 543
rect 19048 757 19082 791
rect 18452 633 18486 667
rect 17800 509 17834 543
rect 21544 757 21578 791
rect 20948 633 20982 667
rect 20296 509 20330 543
rect 2228 385 2262 419
rect 4724 385 4758 419
rect 7220 385 7254 419
rect 9716 385 9750 419
rect 12212 385 12246 419
rect 14708 385 14742 419
rect 17204 385 17238 419
rect 19700 385 19734 419
<< locali >>
rect 4072 791 4106 807
rect 4072 741 4106 757
rect 6568 791 6602 807
rect 6568 741 6602 757
rect 9064 791 9098 807
rect 9064 741 9098 757
rect 11560 791 11594 807
rect 11560 741 11594 757
rect 14056 791 14090 807
rect 14056 741 14090 757
rect 16552 791 16586 807
rect 16552 741 16586 757
rect 19048 791 19082 807
rect 19048 741 19082 757
rect 21544 791 21578 807
rect 21544 741 21578 757
rect 3476 667 3510 683
rect 3476 617 3510 633
rect 5972 667 6006 683
rect 5972 617 6006 633
rect 8468 667 8502 683
rect 8468 617 8502 633
rect 10964 667 10998 683
rect 10964 617 10998 633
rect 13460 667 13494 683
rect 13460 617 13494 633
rect 15956 667 15990 683
rect 15956 617 15990 633
rect 18452 667 18486 683
rect 18452 617 18486 633
rect 20948 667 20982 683
rect 20948 617 20982 633
rect 2824 543 2858 559
rect 2824 493 2858 509
rect 5320 543 5354 559
rect 5320 493 5354 509
rect 7816 543 7850 559
rect 7816 493 7850 509
rect 10312 543 10346 559
rect 10312 493 10346 509
rect 12808 543 12842 559
rect 12808 493 12842 509
rect 15304 543 15338 559
rect 15304 493 15338 509
rect 17800 543 17834 559
rect 17800 493 17834 509
rect 20296 543 20330 559
rect 20296 493 20330 509
rect 2228 419 2262 435
rect 2228 369 2262 385
rect 4724 419 4758 435
rect 4724 369 4758 385
rect 7220 419 7254 435
rect 7220 369 7254 385
rect 9716 419 9750 435
rect 9716 369 9750 385
rect 12212 419 12246 435
rect 12212 369 12246 385
rect 14708 419 14742 435
rect 14708 369 14742 385
rect 17204 419 17238 435
rect 17204 369 17238 385
rect 19700 419 19734 435
rect 19700 369 19734 385
<< viali >>
rect 4072 757 4106 791
rect 6568 757 6602 791
rect 9064 757 9098 791
rect 11560 757 11594 791
rect 14056 757 14090 791
rect 16552 757 16586 791
rect 19048 757 19082 791
rect 21544 757 21578 791
rect 3476 633 3510 667
rect 5972 633 6006 667
rect 8468 633 8502 667
rect 10964 633 10998 667
rect 13460 633 13494 667
rect 15956 633 15990 667
rect 18452 633 18486 667
rect 20948 633 20982 667
rect 2824 509 2858 543
rect 5320 509 5354 543
rect 7816 509 7850 543
rect 10312 509 10346 543
rect 12808 509 12842 543
rect 15304 509 15338 543
rect 17800 509 17834 543
rect 20296 509 20330 543
rect 2228 385 2262 419
rect 4724 385 4758 419
rect 7220 385 7254 419
rect 9716 385 9750 419
rect 12212 385 12246 419
rect 14708 385 14742 419
rect 17204 385 17238 419
rect 19700 385 19734 419
<< metal1 >>
rect 1999 2128 2027 2184
rect 2463 2128 2491 2184
rect 2595 2128 2623 2184
rect 3059 2128 3087 2184
rect 3247 2128 3275 2184
rect 3711 2128 3739 2184
rect 3843 2128 3871 2184
rect 4307 2128 4335 2184
rect 4495 2128 4523 2184
rect 4959 2128 4987 2184
rect 5091 2128 5119 2184
rect 5555 2128 5583 2184
rect 5743 2128 5771 2184
rect 6207 2128 6235 2184
rect 6339 2128 6367 2184
rect 6803 2128 6831 2184
rect 6991 2128 7019 2184
rect 7455 2128 7483 2184
rect 7587 2128 7615 2184
rect 8051 2128 8079 2184
rect 8239 2128 8267 2184
rect 8703 2128 8731 2184
rect 8835 2128 8863 2184
rect 9299 2128 9327 2184
rect 9487 2128 9515 2184
rect 9951 2128 9979 2184
rect 10083 2128 10111 2184
rect 10547 2128 10575 2184
rect 10735 2128 10763 2184
rect 11199 2128 11227 2184
rect 11331 2128 11359 2184
rect 11795 2128 11823 2184
rect 11983 2128 12011 2184
rect 12447 2128 12475 2184
rect 12579 2128 12607 2184
rect 13043 2128 13071 2184
rect 13231 2128 13259 2184
rect 13695 2128 13723 2184
rect 13827 2128 13855 2184
rect 14291 2128 14319 2184
rect 14479 2128 14507 2184
rect 14943 2128 14971 2184
rect 15075 2128 15103 2184
rect 15539 2128 15567 2184
rect 15727 2128 15755 2184
rect 16191 2128 16219 2184
rect 16323 2128 16351 2184
rect 16787 2128 16815 2184
rect 16975 2128 17003 2184
rect 17439 2128 17467 2184
rect 17571 2128 17599 2184
rect 18035 2128 18063 2184
rect 18223 2128 18251 2184
rect 18687 2128 18715 2184
rect 18819 2128 18847 2184
rect 19283 2128 19311 2184
rect 19471 2128 19499 2184
rect 19935 2128 19963 2184
rect 20067 2128 20095 2184
rect 20531 2128 20559 2184
rect 20719 2128 20747 2184
rect 21183 2128 21211 2184
rect 21315 2128 21343 2184
rect 21779 2128 21807 2184
rect 2511 1505 2517 1557
rect 2569 1505 2575 1557
rect 3759 1505 3765 1557
rect 3817 1505 3823 1557
rect 5007 1505 5013 1557
rect 5065 1505 5071 1557
rect 6255 1505 6261 1557
rect 6313 1505 6319 1557
rect 7503 1505 7509 1557
rect 7561 1505 7567 1557
rect 8751 1505 8757 1557
rect 8809 1505 8815 1557
rect 9999 1505 10005 1557
rect 10057 1505 10063 1557
rect 11247 1505 11253 1557
rect 11305 1505 11311 1557
rect 12495 1505 12501 1557
rect 12553 1505 12559 1557
rect 13743 1505 13749 1557
rect 13801 1505 13807 1557
rect 14991 1505 14997 1557
rect 15049 1505 15055 1557
rect 16239 1505 16245 1557
rect 16297 1505 16303 1557
rect 17487 1505 17493 1557
rect 17545 1505 17551 1557
rect 18735 1505 18741 1557
rect 18793 1505 18799 1557
rect 19983 1505 19989 1557
rect 20041 1505 20047 1557
rect 21231 1505 21237 1557
rect 21289 1505 21295 1557
rect 1999 274 2027 868
rect 2213 376 2219 428
rect 2271 376 2277 428
rect 1981 222 1987 274
rect 2039 222 2045 274
rect 2463 150 2491 868
rect 2595 150 2623 868
rect 2809 500 2815 552
rect 2867 500 2873 552
rect 3059 274 3087 868
rect 3247 274 3275 868
rect 3461 624 3467 676
rect 3519 624 3525 676
rect 3041 222 3047 274
rect 3099 222 3105 274
rect 3229 222 3235 274
rect 3287 222 3293 274
rect 3711 150 3739 868
rect 3843 150 3871 868
rect 4057 748 4063 800
rect 4115 748 4121 800
rect 4307 274 4335 868
rect 4495 274 4523 868
rect 4709 376 4715 428
rect 4767 376 4773 428
rect 4289 222 4295 274
rect 4347 222 4353 274
rect 4477 222 4483 274
rect 4535 222 4541 274
rect 4959 150 4987 868
rect 5091 150 5119 868
rect 5305 500 5311 552
rect 5363 500 5369 552
rect 5555 274 5583 868
rect 5743 274 5771 868
rect 5957 624 5963 676
rect 6015 624 6021 676
rect 5537 222 5543 274
rect 5595 222 5601 274
rect 5725 222 5731 274
rect 5783 222 5789 274
rect 6207 150 6235 868
rect 6339 150 6367 868
rect 6553 748 6559 800
rect 6611 748 6617 800
rect 6803 274 6831 868
rect 6991 274 7019 868
rect 7205 376 7211 428
rect 7263 376 7269 428
rect 6785 222 6791 274
rect 6843 222 6849 274
rect 6973 222 6979 274
rect 7031 222 7037 274
rect 7455 150 7483 868
rect 7587 150 7615 868
rect 7801 500 7807 552
rect 7859 500 7865 552
rect 8051 274 8079 868
rect 8239 274 8267 868
rect 8453 624 8459 676
rect 8511 624 8517 676
rect 8033 222 8039 274
rect 8091 222 8097 274
rect 8221 222 8227 274
rect 8279 222 8285 274
rect 8703 150 8731 868
rect 8835 150 8863 868
rect 9049 748 9055 800
rect 9107 748 9113 800
rect 9299 274 9327 868
rect 9487 274 9515 868
rect 9701 376 9707 428
rect 9759 376 9765 428
rect 9281 222 9287 274
rect 9339 222 9345 274
rect 9469 222 9475 274
rect 9527 222 9533 274
rect 9951 150 9979 868
rect 10083 150 10111 868
rect 10297 500 10303 552
rect 10355 500 10361 552
rect 10547 274 10575 868
rect 10735 274 10763 868
rect 10949 624 10955 676
rect 11007 624 11013 676
rect 10529 222 10535 274
rect 10587 222 10593 274
rect 10717 222 10723 274
rect 10775 222 10781 274
rect 11199 150 11227 868
rect 11331 150 11359 868
rect 11545 748 11551 800
rect 11603 748 11609 800
rect 11795 274 11823 868
rect 11983 274 12011 868
rect 12197 376 12203 428
rect 12255 376 12261 428
rect 11777 222 11783 274
rect 11835 222 11841 274
rect 11965 222 11971 274
rect 12023 222 12029 274
rect 12447 150 12475 868
rect 12579 150 12607 868
rect 12793 500 12799 552
rect 12851 500 12857 552
rect 13043 274 13071 868
rect 13231 274 13259 868
rect 13445 624 13451 676
rect 13503 624 13509 676
rect 13025 222 13031 274
rect 13083 222 13089 274
rect 13213 222 13219 274
rect 13271 222 13277 274
rect 13695 150 13723 868
rect 13827 150 13855 868
rect 14041 748 14047 800
rect 14099 748 14105 800
rect 14291 274 14319 868
rect 14479 274 14507 868
rect 14693 376 14699 428
rect 14751 376 14757 428
rect 14273 222 14279 274
rect 14331 222 14337 274
rect 14461 222 14467 274
rect 14519 222 14525 274
rect 14943 150 14971 868
rect 15075 150 15103 868
rect 15289 500 15295 552
rect 15347 500 15353 552
rect 15539 274 15567 868
rect 15727 274 15755 868
rect 15941 624 15947 676
rect 15999 624 16005 676
rect 15521 222 15527 274
rect 15579 222 15585 274
rect 15709 222 15715 274
rect 15767 222 15773 274
rect 16191 150 16219 868
rect 16323 150 16351 868
rect 16537 748 16543 800
rect 16595 748 16601 800
rect 16787 274 16815 868
rect 16975 274 17003 868
rect 17189 376 17195 428
rect 17247 376 17253 428
rect 16769 222 16775 274
rect 16827 222 16833 274
rect 16957 222 16963 274
rect 17015 222 17021 274
rect 17439 150 17467 868
rect 17571 150 17599 868
rect 17785 500 17791 552
rect 17843 500 17849 552
rect 18035 274 18063 868
rect 18223 274 18251 868
rect 18437 624 18443 676
rect 18495 624 18501 676
rect 18017 222 18023 274
rect 18075 222 18081 274
rect 18205 222 18211 274
rect 18263 222 18269 274
rect 18687 150 18715 868
rect 18819 150 18847 868
rect 19033 748 19039 800
rect 19091 748 19097 800
rect 19283 274 19311 868
rect 19471 274 19499 868
rect 19685 376 19691 428
rect 19743 376 19749 428
rect 19265 222 19271 274
rect 19323 222 19329 274
rect 19453 222 19459 274
rect 19511 222 19517 274
rect 19935 150 19963 868
rect 20067 150 20095 868
rect 20281 500 20287 552
rect 20339 500 20345 552
rect 20531 274 20559 868
rect 20719 274 20747 868
rect 20933 624 20939 676
rect 20991 624 20997 676
rect 20513 222 20519 274
rect 20571 222 20577 274
rect 20701 222 20707 274
rect 20759 222 20765 274
rect 21183 150 21211 868
rect 21315 150 21343 868
rect 21529 748 21535 800
rect 21587 748 21593 800
rect 21779 274 21807 868
rect 21761 222 21767 274
rect 21819 222 21825 274
rect 2445 98 2451 150
rect 2503 98 2509 150
rect 2577 98 2583 150
rect 2635 98 2641 150
rect 3693 98 3699 150
rect 3751 98 3757 150
rect 3825 98 3831 150
rect 3883 98 3889 150
rect 4941 98 4947 150
rect 4999 98 5005 150
rect 5073 98 5079 150
rect 5131 98 5137 150
rect 6189 98 6195 150
rect 6247 98 6253 150
rect 6321 98 6327 150
rect 6379 98 6385 150
rect 7437 98 7443 150
rect 7495 98 7501 150
rect 7569 98 7575 150
rect 7627 98 7633 150
rect 8685 98 8691 150
rect 8743 98 8749 150
rect 8817 98 8823 150
rect 8875 98 8881 150
rect 9933 98 9939 150
rect 9991 98 9997 150
rect 10065 98 10071 150
rect 10123 98 10129 150
rect 11181 98 11187 150
rect 11239 98 11245 150
rect 11313 98 11319 150
rect 11371 98 11377 150
rect 12429 98 12435 150
rect 12487 98 12493 150
rect 12561 98 12567 150
rect 12619 98 12625 150
rect 13677 98 13683 150
rect 13735 98 13741 150
rect 13809 98 13815 150
rect 13867 98 13873 150
rect 14925 98 14931 150
rect 14983 98 14989 150
rect 15057 98 15063 150
rect 15115 98 15121 150
rect 16173 98 16179 150
rect 16231 98 16237 150
rect 16305 98 16311 150
rect 16363 98 16369 150
rect 17421 98 17427 150
rect 17479 98 17485 150
rect 17553 98 17559 150
rect 17611 98 17617 150
rect 18669 98 18675 150
rect 18727 98 18733 150
rect 18801 98 18807 150
rect 18859 98 18865 150
rect 19917 98 19923 150
rect 19975 98 19981 150
rect 20049 98 20055 150
rect 20107 98 20113 150
rect 21165 98 21171 150
rect 21223 98 21229 150
rect 21297 98 21303 150
rect 21355 98 21361 150
<< via1 >>
rect 2517 1505 2569 1557
rect 3765 1505 3817 1557
rect 5013 1505 5065 1557
rect 6261 1505 6313 1557
rect 7509 1505 7561 1557
rect 8757 1505 8809 1557
rect 10005 1505 10057 1557
rect 11253 1505 11305 1557
rect 12501 1505 12553 1557
rect 13749 1505 13801 1557
rect 14997 1505 15049 1557
rect 16245 1505 16297 1557
rect 17493 1505 17545 1557
rect 18741 1505 18793 1557
rect 19989 1505 20041 1557
rect 21237 1505 21289 1557
rect 2219 419 2271 428
rect 2219 385 2228 419
rect 2228 385 2262 419
rect 2262 385 2271 419
rect 2219 376 2271 385
rect 1987 222 2039 274
rect 2815 543 2867 552
rect 2815 509 2824 543
rect 2824 509 2858 543
rect 2858 509 2867 543
rect 2815 500 2867 509
rect 3467 667 3519 676
rect 3467 633 3476 667
rect 3476 633 3510 667
rect 3510 633 3519 667
rect 3467 624 3519 633
rect 3047 222 3099 274
rect 3235 222 3287 274
rect 4063 791 4115 800
rect 4063 757 4072 791
rect 4072 757 4106 791
rect 4106 757 4115 791
rect 4063 748 4115 757
rect 4715 419 4767 428
rect 4715 385 4724 419
rect 4724 385 4758 419
rect 4758 385 4767 419
rect 4715 376 4767 385
rect 4295 222 4347 274
rect 4483 222 4535 274
rect 5311 543 5363 552
rect 5311 509 5320 543
rect 5320 509 5354 543
rect 5354 509 5363 543
rect 5311 500 5363 509
rect 5963 667 6015 676
rect 5963 633 5972 667
rect 5972 633 6006 667
rect 6006 633 6015 667
rect 5963 624 6015 633
rect 5543 222 5595 274
rect 5731 222 5783 274
rect 6559 791 6611 800
rect 6559 757 6568 791
rect 6568 757 6602 791
rect 6602 757 6611 791
rect 6559 748 6611 757
rect 7211 419 7263 428
rect 7211 385 7220 419
rect 7220 385 7254 419
rect 7254 385 7263 419
rect 7211 376 7263 385
rect 6791 222 6843 274
rect 6979 222 7031 274
rect 7807 543 7859 552
rect 7807 509 7816 543
rect 7816 509 7850 543
rect 7850 509 7859 543
rect 7807 500 7859 509
rect 8459 667 8511 676
rect 8459 633 8468 667
rect 8468 633 8502 667
rect 8502 633 8511 667
rect 8459 624 8511 633
rect 8039 222 8091 274
rect 8227 222 8279 274
rect 9055 791 9107 800
rect 9055 757 9064 791
rect 9064 757 9098 791
rect 9098 757 9107 791
rect 9055 748 9107 757
rect 9707 419 9759 428
rect 9707 385 9716 419
rect 9716 385 9750 419
rect 9750 385 9759 419
rect 9707 376 9759 385
rect 9287 222 9339 274
rect 9475 222 9527 274
rect 10303 543 10355 552
rect 10303 509 10312 543
rect 10312 509 10346 543
rect 10346 509 10355 543
rect 10303 500 10355 509
rect 10955 667 11007 676
rect 10955 633 10964 667
rect 10964 633 10998 667
rect 10998 633 11007 667
rect 10955 624 11007 633
rect 10535 222 10587 274
rect 10723 222 10775 274
rect 11551 791 11603 800
rect 11551 757 11560 791
rect 11560 757 11594 791
rect 11594 757 11603 791
rect 11551 748 11603 757
rect 12203 419 12255 428
rect 12203 385 12212 419
rect 12212 385 12246 419
rect 12246 385 12255 419
rect 12203 376 12255 385
rect 11783 222 11835 274
rect 11971 222 12023 274
rect 12799 543 12851 552
rect 12799 509 12808 543
rect 12808 509 12842 543
rect 12842 509 12851 543
rect 12799 500 12851 509
rect 13451 667 13503 676
rect 13451 633 13460 667
rect 13460 633 13494 667
rect 13494 633 13503 667
rect 13451 624 13503 633
rect 13031 222 13083 274
rect 13219 222 13271 274
rect 14047 791 14099 800
rect 14047 757 14056 791
rect 14056 757 14090 791
rect 14090 757 14099 791
rect 14047 748 14099 757
rect 14699 419 14751 428
rect 14699 385 14708 419
rect 14708 385 14742 419
rect 14742 385 14751 419
rect 14699 376 14751 385
rect 14279 222 14331 274
rect 14467 222 14519 274
rect 15295 543 15347 552
rect 15295 509 15304 543
rect 15304 509 15338 543
rect 15338 509 15347 543
rect 15295 500 15347 509
rect 15947 667 15999 676
rect 15947 633 15956 667
rect 15956 633 15990 667
rect 15990 633 15999 667
rect 15947 624 15999 633
rect 15527 222 15579 274
rect 15715 222 15767 274
rect 16543 791 16595 800
rect 16543 757 16552 791
rect 16552 757 16586 791
rect 16586 757 16595 791
rect 16543 748 16595 757
rect 17195 419 17247 428
rect 17195 385 17204 419
rect 17204 385 17238 419
rect 17238 385 17247 419
rect 17195 376 17247 385
rect 16775 222 16827 274
rect 16963 222 17015 274
rect 17791 543 17843 552
rect 17791 509 17800 543
rect 17800 509 17834 543
rect 17834 509 17843 543
rect 17791 500 17843 509
rect 18443 667 18495 676
rect 18443 633 18452 667
rect 18452 633 18486 667
rect 18486 633 18495 667
rect 18443 624 18495 633
rect 18023 222 18075 274
rect 18211 222 18263 274
rect 19039 791 19091 800
rect 19039 757 19048 791
rect 19048 757 19082 791
rect 19082 757 19091 791
rect 19039 748 19091 757
rect 19691 419 19743 428
rect 19691 385 19700 419
rect 19700 385 19734 419
rect 19734 385 19743 419
rect 19691 376 19743 385
rect 19271 222 19323 274
rect 19459 222 19511 274
rect 20287 543 20339 552
rect 20287 509 20296 543
rect 20296 509 20330 543
rect 20330 509 20339 543
rect 20287 500 20339 509
rect 20939 667 20991 676
rect 20939 633 20948 667
rect 20948 633 20982 667
rect 20982 633 20991 667
rect 20939 624 20991 633
rect 20519 222 20571 274
rect 20707 222 20759 274
rect 21535 791 21587 800
rect 21535 757 21544 791
rect 21544 757 21578 791
rect 21578 757 21587 791
rect 21535 748 21587 757
rect 21767 222 21819 274
rect 2451 98 2503 150
rect 2583 98 2635 150
rect 3699 98 3751 150
rect 3831 98 3883 150
rect 4947 98 4999 150
rect 5079 98 5131 150
rect 6195 98 6247 150
rect 6327 98 6379 150
rect 7443 98 7495 150
rect 7575 98 7627 150
rect 8691 98 8743 150
rect 8823 98 8875 150
rect 9939 98 9991 150
rect 10071 98 10123 150
rect 11187 98 11239 150
rect 11319 98 11371 150
rect 12435 98 12487 150
rect 12567 98 12619 150
rect 13683 98 13735 150
rect 13815 98 13867 150
rect 14931 98 14983 150
rect 15063 98 15115 150
rect 16179 98 16231 150
rect 16311 98 16363 150
rect 17427 98 17479 150
rect 17559 98 17611 150
rect 18675 98 18727 150
rect 18807 98 18859 150
rect 19923 98 19975 150
rect 20055 98 20107 150
rect 21171 98 21223 150
rect 21303 98 21355 150
<< metal2 >>
rect 2515 1559 2571 1568
rect 2515 1494 2571 1503
rect 3763 1559 3819 1568
rect 3763 1494 3819 1503
rect 5011 1559 5067 1568
rect 5011 1494 5067 1503
rect 6259 1559 6315 1568
rect 6259 1494 6315 1503
rect 7507 1559 7563 1568
rect 7507 1494 7563 1503
rect 8755 1559 8811 1568
rect 8755 1494 8811 1503
rect 10003 1559 10059 1568
rect 10003 1494 10059 1503
rect 11251 1559 11307 1568
rect 11251 1494 11307 1503
rect 12499 1559 12555 1568
rect 12499 1494 12555 1503
rect 13747 1559 13803 1568
rect 13747 1494 13803 1503
rect 14995 1559 15051 1568
rect 14995 1494 15051 1503
rect 16243 1559 16299 1568
rect 16243 1494 16299 1503
rect 17491 1559 17547 1568
rect 17491 1494 17547 1503
rect 18739 1559 18795 1568
rect 18739 1494 18795 1503
rect 19987 1559 20043 1568
rect 19987 1494 20043 1503
rect 21235 1559 21291 1568
rect 21235 1494 21291 1503
rect 4061 802 4117 811
rect 4061 737 4117 746
rect 6557 802 6613 811
rect 6557 737 6613 746
rect 9053 802 9109 811
rect 9053 737 9109 746
rect 11549 802 11605 811
rect 11549 737 11605 746
rect 14045 802 14101 811
rect 14045 737 14101 746
rect 16541 802 16597 811
rect 16541 737 16597 746
rect 19037 802 19093 811
rect 19037 737 19093 746
rect 21533 802 21589 811
rect 21533 737 21589 746
rect 3465 678 3521 687
rect 3465 613 3521 622
rect 5961 678 6017 687
rect 5961 613 6017 622
rect 8457 678 8513 687
rect 8457 613 8513 622
rect 10953 678 11009 687
rect 10953 613 11009 622
rect 13449 678 13505 687
rect 13449 613 13505 622
rect 15945 678 16001 687
rect 15945 613 16001 622
rect 18441 678 18497 687
rect 18441 613 18497 622
rect 20937 678 20993 687
rect 20937 613 20993 622
rect 2813 554 2869 563
rect 2813 489 2869 498
rect 5309 554 5365 563
rect 5309 489 5365 498
rect 7805 554 7861 563
rect 7805 489 7861 498
rect 10301 554 10357 563
rect 10301 489 10357 498
rect 12797 554 12853 563
rect 12797 489 12853 498
rect 15293 554 15349 563
rect 15293 489 15349 498
rect 17789 554 17845 563
rect 17789 489 17845 498
rect 20285 554 20341 563
rect 20285 489 20341 498
rect 2217 430 2273 439
rect 2217 365 2273 374
rect 4713 430 4769 439
rect 4713 365 4769 374
rect 7209 430 7265 439
rect 7209 365 7265 374
rect 9705 430 9761 439
rect 9705 365 9761 374
rect 12201 430 12257 439
rect 12201 365 12257 374
rect 14697 430 14753 439
rect 14697 365 14753 374
rect 17193 430 17249 439
rect 17193 365 17249 374
rect 19689 430 19745 439
rect 19689 365 19745 374
rect 1985 276 2041 285
rect 1985 211 2041 220
rect 3045 276 3101 285
rect 3045 211 3101 220
rect 3233 276 3289 285
rect 3233 211 3289 220
rect 4293 276 4349 285
rect 4293 211 4349 220
rect 4481 276 4537 285
rect 4481 211 4537 220
rect 5541 276 5597 285
rect 5541 211 5597 220
rect 5729 276 5785 285
rect 5729 211 5785 220
rect 6789 276 6845 285
rect 6789 211 6845 220
rect 6977 276 7033 285
rect 6977 211 7033 220
rect 8037 276 8093 285
rect 8037 211 8093 220
rect 8225 276 8281 285
rect 8225 211 8281 220
rect 9285 276 9341 285
rect 9285 211 9341 220
rect 9473 276 9529 285
rect 9473 211 9529 220
rect 10533 276 10589 285
rect 10533 211 10589 220
rect 10721 276 10777 285
rect 10721 211 10777 220
rect 11781 276 11837 285
rect 11781 211 11837 220
rect 11969 276 12025 285
rect 11969 211 12025 220
rect 13029 276 13085 285
rect 13029 211 13085 220
rect 13217 276 13273 285
rect 13217 211 13273 220
rect 14277 276 14333 285
rect 14277 211 14333 220
rect 14465 276 14521 285
rect 14465 211 14521 220
rect 15525 276 15581 285
rect 15525 211 15581 220
rect 15713 276 15769 285
rect 15713 211 15769 220
rect 16773 276 16829 285
rect 16773 211 16829 220
rect 16961 276 17017 285
rect 16961 211 17017 220
rect 18021 276 18077 285
rect 18021 211 18077 220
rect 18209 276 18265 285
rect 18209 211 18265 220
rect 19269 276 19325 285
rect 19269 211 19325 220
rect 19457 276 19513 285
rect 19457 211 19513 220
rect 20517 276 20573 285
rect 20517 211 20573 220
rect 20705 276 20761 285
rect 20705 211 20761 220
rect 21765 276 21821 285
rect 21765 211 21821 220
rect 2449 152 2505 161
rect 2449 87 2505 96
rect 2581 152 2637 161
rect 2581 87 2637 96
rect 3697 152 3753 161
rect 3697 87 3753 96
rect 3829 152 3885 161
rect 3829 87 3885 96
rect 4945 152 5001 161
rect 4945 87 5001 96
rect 5077 152 5133 161
rect 5077 87 5133 96
rect 6193 152 6249 161
rect 6193 87 6249 96
rect 6325 152 6381 161
rect 6325 87 6381 96
rect 7441 152 7497 161
rect 7441 87 7497 96
rect 7573 152 7629 161
rect 7573 87 7629 96
rect 8689 152 8745 161
rect 8689 87 8745 96
rect 8821 152 8877 161
rect 8821 87 8877 96
rect 9937 152 9993 161
rect 9937 87 9993 96
rect 10069 152 10125 161
rect 10069 87 10125 96
rect 11185 152 11241 161
rect 11185 87 11241 96
rect 11317 152 11373 161
rect 11317 87 11373 96
rect 12433 152 12489 161
rect 12433 87 12489 96
rect 12565 152 12621 161
rect 12565 87 12621 96
rect 13681 152 13737 161
rect 13681 87 13737 96
rect 13813 152 13869 161
rect 13813 87 13869 96
rect 14929 152 14985 161
rect 14929 87 14985 96
rect 15061 152 15117 161
rect 15061 87 15117 96
rect 16177 152 16233 161
rect 16177 87 16233 96
rect 16309 152 16365 161
rect 16309 87 16365 96
rect 17425 152 17481 161
rect 17425 87 17481 96
rect 17557 152 17613 161
rect 17557 87 17613 96
rect 18673 152 18729 161
rect 18673 87 18729 96
rect 18805 152 18861 161
rect 18805 87 18861 96
rect 19921 152 19977 161
rect 19921 87 19977 96
rect 20053 152 20109 161
rect 20053 87 20109 96
rect 21169 152 21225 161
rect 21169 87 21225 96
rect 21301 152 21357 161
rect 21301 87 21357 96
<< via2 >>
rect 2515 1557 2571 1559
rect 2515 1505 2517 1557
rect 2517 1505 2569 1557
rect 2569 1505 2571 1557
rect 2515 1503 2571 1505
rect 3763 1557 3819 1559
rect 3763 1505 3765 1557
rect 3765 1505 3817 1557
rect 3817 1505 3819 1557
rect 3763 1503 3819 1505
rect 5011 1557 5067 1559
rect 5011 1505 5013 1557
rect 5013 1505 5065 1557
rect 5065 1505 5067 1557
rect 5011 1503 5067 1505
rect 6259 1557 6315 1559
rect 6259 1505 6261 1557
rect 6261 1505 6313 1557
rect 6313 1505 6315 1557
rect 6259 1503 6315 1505
rect 7507 1557 7563 1559
rect 7507 1505 7509 1557
rect 7509 1505 7561 1557
rect 7561 1505 7563 1557
rect 7507 1503 7563 1505
rect 8755 1557 8811 1559
rect 8755 1505 8757 1557
rect 8757 1505 8809 1557
rect 8809 1505 8811 1557
rect 8755 1503 8811 1505
rect 10003 1557 10059 1559
rect 10003 1505 10005 1557
rect 10005 1505 10057 1557
rect 10057 1505 10059 1557
rect 10003 1503 10059 1505
rect 11251 1557 11307 1559
rect 11251 1505 11253 1557
rect 11253 1505 11305 1557
rect 11305 1505 11307 1557
rect 11251 1503 11307 1505
rect 12499 1557 12555 1559
rect 12499 1505 12501 1557
rect 12501 1505 12553 1557
rect 12553 1505 12555 1557
rect 12499 1503 12555 1505
rect 13747 1557 13803 1559
rect 13747 1505 13749 1557
rect 13749 1505 13801 1557
rect 13801 1505 13803 1557
rect 13747 1503 13803 1505
rect 14995 1557 15051 1559
rect 14995 1505 14997 1557
rect 14997 1505 15049 1557
rect 15049 1505 15051 1557
rect 14995 1503 15051 1505
rect 16243 1557 16299 1559
rect 16243 1505 16245 1557
rect 16245 1505 16297 1557
rect 16297 1505 16299 1557
rect 16243 1503 16299 1505
rect 17491 1557 17547 1559
rect 17491 1505 17493 1557
rect 17493 1505 17545 1557
rect 17545 1505 17547 1557
rect 17491 1503 17547 1505
rect 18739 1557 18795 1559
rect 18739 1505 18741 1557
rect 18741 1505 18793 1557
rect 18793 1505 18795 1557
rect 18739 1503 18795 1505
rect 19987 1557 20043 1559
rect 19987 1505 19989 1557
rect 19989 1505 20041 1557
rect 20041 1505 20043 1557
rect 19987 1503 20043 1505
rect 21235 1557 21291 1559
rect 21235 1505 21237 1557
rect 21237 1505 21289 1557
rect 21289 1505 21291 1557
rect 21235 1503 21291 1505
rect 4061 800 4117 802
rect 4061 748 4063 800
rect 4063 748 4115 800
rect 4115 748 4117 800
rect 4061 746 4117 748
rect 6557 800 6613 802
rect 6557 748 6559 800
rect 6559 748 6611 800
rect 6611 748 6613 800
rect 6557 746 6613 748
rect 9053 800 9109 802
rect 9053 748 9055 800
rect 9055 748 9107 800
rect 9107 748 9109 800
rect 9053 746 9109 748
rect 11549 800 11605 802
rect 11549 748 11551 800
rect 11551 748 11603 800
rect 11603 748 11605 800
rect 11549 746 11605 748
rect 14045 800 14101 802
rect 14045 748 14047 800
rect 14047 748 14099 800
rect 14099 748 14101 800
rect 14045 746 14101 748
rect 16541 800 16597 802
rect 16541 748 16543 800
rect 16543 748 16595 800
rect 16595 748 16597 800
rect 16541 746 16597 748
rect 19037 800 19093 802
rect 19037 748 19039 800
rect 19039 748 19091 800
rect 19091 748 19093 800
rect 19037 746 19093 748
rect 21533 800 21589 802
rect 21533 748 21535 800
rect 21535 748 21587 800
rect 21587 748 21589 800
rect 21533 746 21589 748
rect 3465 676 3521 678
rect 3465 624 3467 676
rect 3467 624 3519 676
rect 3519 624 3521 676
rect 3465 622 3521 624
rect 5961 676 6017 678
rect 5961 624 5963 676
rect 5963 624 6015 676
rect 6015 624 6017 676
rect 5961 622 6017 624
rect 8457 676 8513 678
rect 8457 624 8459 676
rect 8459 624 8511 676
rect 8511 624 8513 676
rect 8457 622 8513 624
rect 10953 676 11009 678
rect 10953 624 10955 676
rect 10955 624 11007 676
rect 11007 624 11009 676
rect 10953 622 11009 624
rect 13449 676 13505 678
rect 13449 624 13451 676
rect 13451 624 13503 676
rect 13503 624 13505 676
rect 13449 622 13505 624
rect 15945 676 16001 678
rect 15945 624 15947 676
rect 15947 624 15999 676
rect 15999 624 16001 676
rect 15945 622 16001 624
rect 18441 676 18497 678
rect 18441 624 18443 676
rect 18443 624 18495 676
rect 18495 624 18497 676
rect 18441 622 18497 624
rect 20937 676 20993 678
rect 20937 624 20939 676
rect 20939 624 20991 676
rect 20991 624 20993 676
rect 20937 622 20993 624
rect 2813 552 2869 554
rect 2813 500 2815 552
rect 2815 500 2867 552
rect 2867 500 2869 552
rect 2813 498 2869 500
rect 5309 552 5365 554
rect 5309 500 5311 552
rect 5311 500 5363 552
rect 5363 500 5365 552
rect 5309 498 5365 500
rect 7805 552 7861 554
rect 7805 500 7807 552
rect 7807 500 7859 552
rect 7859 500 7861 552
rect 7805 498 7861 500
rect 10301 552 10357 554
rect 10301 500 10303 552
rect 10303 500 10355 552
rect 10355 500 10357 552
rect 10301 498 10357 500
rect 12797 552 12853 554
rect 12797 500 12799 552
rect 12799 500 12851 552
rect 12851 500 12853 552
rect 12797 498 12853 500
rect 15293 552 15349 554
rect 15293 500 15295 552
rect 15295 500 15347 552
rect 15347 500 15349 552
rect 15293 498 15349 500
rect 17789 552 17845 554
rect 17789 500 17791 552
rect 17791 500 17843 552
rect 17843 500 17845 552
rect 17789 498 17845 500
rect 20285 552 20341 554
rect 20285 500 20287 552
rect 20287 500 20339 552
rect 20339 500 20341 552
rect 20285 498 20341 500
rect 2217 428 2273 430
rect 2217 376 2219 428
rect 2219 376 2271 428
rect 2271 376 2273 428
rect 2217 374 2273 376
rect 4713 428 4769 430
rect 4713 376 4715 428
rect 4715 376 4767 428
rect 4767 376 4769 428
rect 4713 374 4769 376
rect 7209 428 7265 430
rect 7209 376 7211 428
rect 7211 376 7263 428
rect 7263 376 7265 428
rect 7209 374 7265 376
rect 9705 428 9761 430
rect 9705 376 9707 428
rect 9707 376 9759 428
rect 9759 376 9761 428
rect 9705 374 9761 376
rect 12201 428 12257 430
rect 12201 376 12203 428
rect 12203 376 12255 428
rect 12255 376 12257 428
rect 12201 374 12257 376
rect 14697 428 14753 430
rect 14697 376 14699 428
rect 14699 376 14751 428
rect 14751 376 14753 428
rect 14697 374 14753 376
rect 17193 428 17249 430
rect 17193 376 17195 428
rect 17195 376 17247 428
rect 17247 376 17249 428
rect 17193 374 17249 376
rect 19689 428 19745 430
rect 19689 376 19691 428
rect 19691 376 19743 428
rect 19743 376 19745 428
rect 19689 374 19745 376
rect 1985 274 2041 276
rect 1985 222 1987 274
rect 1987 222 2039 274
rect 2039 222 2041 274
rect 1985 220 2041 222
rect 3045 274 3101 276
rect 3045 222 3047 274
rect 3047 222 3099 274
rect 3099 222 3101 274
rect 3045 220 3101 222
rect 3233 274 3289 276
rect 3233 222 3235 274
rect 3235 222 3287 274
rect 3287 222 3289 274
rect 3233 220 3289 222
rect 4293 274 4349 276
rect 4293 222 4295 274
rect 4295 222 4347 274
rect 4347 222 4349 274
rect 4293 220 4349 222
rect 4481 274 4537 276
rect 4481 222 4483 274
rect 4483 222 4535 274
rect 4535 222 4537 274
rect 4481 220 4537 222
rect 5541 274 5597 276
rect 5541 222 5543 274
rect 5543 222 5595 274
rect 5595 222 5597 274
rect 5541 220 5597 222
rect 5729 274 5785 276
rect 5729 222 5731 274
rect 5731 222 5783 274
rect 5783 222 5785 274
rect 5729 220 5785 222
rect 6789 274 6845 276
rect 6789 222 6791 274
rect 6791 222 6843 274
rect 6843 222 6845 274
rect 6789 220 6845 222
rect 6977 274 7033 276
rect 6977 222 6979 274
rect 6979 222 7031 274
rect 7031 222 7033 274
rect 6977 220 7033 222
rect 8037 274 8093 276
rect 8037 222 8039 274
rect 8039 222 8091 274
rect 8091 222 8093 274
rect 8037 220 8093 222
rect 8225 274 8281 276
rect 8225 222 8227 274
rect 8227 222 8279 274
rect 8279 222 8281 274
rect 8225 220 8281 222
rect 9285 274 9341 276
rect 9285 222 9287 274
rect 9287 222 9339 274
rect 9339 222 9341 274
rect 9285 220 9341 222
rect 9473 274 9529 276
rect 9473 222 9475 274
rect 9475 222 9527 274
rect 9527 222 9529 274
rect 9473 220 9529 222
rect 10533 274 10589 276
rect 10533 222 10535 274
rect 10535 222 10587 274
rect 10587 222 10589 274
rect 10533 220 10589 222
rect 10721 274 10777 276
rect 10721 222 10723 274
rect 10723 222 10775 274
rect 10775 222 10777 274
rect 10721 220 10777 222
rect 11781 274 11837 276
rect 11781 222 11783 274
rect 11783 222 11835 274
rect 11835 222 11837 274
rect 11781 220 11837 222
rect 11969 274 12025 276
rect 11969 222 11971 274
rect 11971 222 12023 274
rect 12023 222 12025 274
rect 11969 220 12025 222
rect 13029 274 13085 276
rect 13029 222 13031 274
rect 13031 222 13083 274
rect 13083 222 13085 274
rect 13029 220 13085 222
rect 13217 274 13273 276
rect 13217 222 13219 274
rect 13219 222 13271 274
rect 13271 222 13273 274
rect 13217 220 13273 222
rect 14277 274 14333 276
rect 14277 222 14279 274
rect 14279 222 14331 274
rect 14331 222 14333 274
rect 14277 220 14333 222
rect 14465 274 14521 276
rect 14465 222 14467 274
rect 14467 222 14519 274
rect 14519 222 14521 274
rect 14465 220 14521 222
rect 15525 274 15581 276
rect 15525 222 15527 274
rect 15527 222 15579 274
rect 15579 222 15581 274
rect 15525 220 15581 222
rect 15713 274 15769 276
rect 15713 222 15715 274
rect 15715 222 15767 274
rect 15767 222 15769 274
rect 15713 220 15769 222
rect 16773 274 16829 276
rect 16773 222 16775 274
rect 16775 222 16827 274
rect 16827 222 16829 274
rect 16773 220 16829 222
rect 16961 274 17017 276
rect 16961 222 16963 274
rect 16963 222 17015 274
rect 17015 222 17017 274
rect 16961 220 17017 222
rect 18021 274 18077 276
rect 18021 222 18023 274
rect 18023 222 18075 274
rect 18075 222 18077 274
rect 18021 220 18077 222
rect 18209 274 18265 276
rect 18209 222 18211 274
rect 18211 222 18263 274
rect 18263 222 18265 274
rect 18209 220 18265 222
rect 19269 274 19325 276
rect 19269 222 19271 274
rect 19271 222 19323 274
rect 19323 222 19325 274
rect 19269 220 19325 222
rect 19457 274 19513 276
rect 19457 222 19459 274
rect 19459 222 19511 274
rect 19511 222 19513 274
rect 19457 220 19513 222
rect 20517 274 20573 276
rect 20517 222 20519 274
rect 20519 222 20571 274
rect 20571 222 20573 274
rect 20517 220 20573 222
rect 20705 274 20761 276
rect 20705 222 20707 274
rect 20707 222 20759 274
rect 20759 222 20761 274
rect 20705 220 20761 222
rect 21765 274 21821 276
rect 21765 222 21767 274
rect 21767 222 21819 274
rect 21819 222 21821 274
rect 21765 220 21821 222
rect 2449 150 2505 152
rect 2449 98 2451 150
rect 2451 98 2503 150
rect 2503 98 2505 150
rect 2449 96 2505 98
rect 2581 150 2637 152
rect 2581 98 2583 150
rect 2583 98 2635 150
rect 2635 98 2637 150
rect 2581 96 2637 98
rect 3697 150 3753 152
rect 3697 98 3699 150
rect 3699 98 3751 150
rect 3751 98 3753 150
rect 3697 96 3753 98
rect 3829 150 3885 152
rect 3829 98 3831 150
rect 3831 98 3883 150
rect 3883 98 3885 150
rect 3829 96 3885 98
rect 4945 150 5001 152
rect 4945 98 4947 150
rect 4947 98 4999 150
rect 4999 98 5001 150
rect 4945 96 5001 98
rect 5077 150 5133 152
rect 5077 98 5079 150
rect 5079 98 5131 150
rect 5131 98 5133 150
rect 5077 96 5133 98
rect 6193 150 6249 152
rect 6193 98 6195 150
rect 6195 98 6247 150
rect 6247 98 6249 150
rect 6193 96 6249 98
rect 6325 150 6381 152
rect 6325 98 6327 150
rect 6327 98 6379 150
rect 6379 98 6381 150
rect 6325 96 6381 98
rect 7441 150 7497 152
rect 7441 98 7443 150
rect 7443 98 7495 150
rect 7495 98 7497 150
rect 7441 96 7497 98
rect 7573 150 7629 152
rect 7573 98 7575 150
rect 7575 98 7627 150
rect 7627 98 7629 150
rect 7573 96 7629 98
rect 8689 150 8745 152
rect 8689 98 8691 150
rect 8691 98 8743 150
rect 8743 98 8745 150
rect 8689 96 8745 98
rect 8821 150 8877 152
rect 8821 98 8823 150
rect 8823 98 8875 150
rect 8875 98 8877 150
rect 8821 96 8877 98
rect 9937 150 9993 152
rect 9937 98 9939 150
rect 9939 98 9991 150
rect 9991 98 9993 150
rect 9937 96 9993 98
rect 10069 150 10125 152
rect 10069 98 10071 150
rect 10071 98 10123 150
rect 10123 98 10125 150
rect 10069 96 10125 98
rect 11185 150 11241 152
rect 11185 98 11187 150
rect 11187 98 11239 150
rect 11239 98 11241 150
rect 11185 96 11241 98
rect 11317 150 11373 152
rect 11317 98 11319 150
rect 11319 98 11371 150
rect 11371 98 11373 150
rect 11317 96 11373 98
rect 12433 150 12489 152
rect 12433 98 12435 150
rect 12435 98 12487 150
rect 12487 98 12489 150
rect 12433 96 12489 98
rect 12565 150 12621 152
rect 12565 98 12567 150
rect 12567 98 12619 150
rect 12619 98 12621 150
rect 12565 96 12621 98
rect 13681 150 13737 152
rect 13681 98 13683 150
rect 13683 98 13735 150
rect 13735 98 13737 150
rect 13681 96 13737 98
rect 13813 150 13869 152
rect 13813 98 13815 150
rect 13815 98 13867 150
rect 13867 98 13869 150
rect 13813 96 13869 98
rect 14929 150 14985 152
rect 14929 98 14931 150
rect 14931 98 14983 150
rect 14983 98 14985 150
rect 14929 96 14985 98
rect 15061 150 15117 152
rect 15061 98 15063 150
rect 15063 98 15115 150
rect 15115 98 15117 150
rect 15061 96 15117 98
rect 16177 150 16233 152
rect 16177 98 16179 150
rect 16179 98 16231 150
rect 16231 98 16233 150
rect 16177 96 16233 98
rect 16309 150 16365 152
rect 16309 98 16311 150
rect 16311 98 16363 150
rect 16363 98 16365 150
rect 16309 96 16365 98
rect 17425 150 17481 152
rect 17425 98 17427 150
rect 17427 98 17479 150
rect 17479 98 17481 150
rect 17425 96 17481 98
rect 17557 150 17613 152
rect 17557 98 17559 150
rect 17559 98 17611 150
rect 17611 98 17613 150
rect 17557 96 17613 98
rect 18673 150 18729 152
rect 18673 98 18675 150
rect 18675 98 18727 150
rect 18727 98 18729 150
rect 18673 96 18729 98
rect 18805 150 18861 152
rect 18805 98 18807 150
rect 18807 98 18859 150
rect 18859 98 18861 150
rect 18805 96 18861 98
rect 19921 150 19977 152
rect 19921 98 19923 150
rect 19923 98 19975 150
rect 19975 98 19977 150
rect 19921 96 19977 98
rect 20053 150 20109 152
rect 20053 98 20055 150
rect 20055 98 20107 150
rect 20107 98 20109 150
rect 20053 96 20109 98
rect 21169 150 21225 152
rect 21169 98 21171 150
rect 21171 98 21223 150
rect 21223 98 21225 150
rect 21169 96 21225 98
rect 21301 150 21357 152
rect 21301 98 21303 150
rect 21303 98 21355 150
rect 21355 98 21357 150
rect 21301 96 21357 98
<< metal3 >>
rect 33 1559 21310 1564
rect 33 1503 2515 1559
rect 2571 1503 3763 1559
rect 3819 1503 5011 1559
rect 5067 1503 6259 1559
rect 6315 1503 7507 1559
rect 7563 1503 8755 1559
rect 8811 1503 10003 1559
rect 10059 1503 11251 1559
rect 11307 1503 12499 1559
rect 12555 1503 13747 1559
rect 13803 1503 14995 1559
rect 15051 1503 16243 1559
rect 16299 1503 17491 1559
rect 17547 1503 18739 1559
rect 18795 1503 19987 1559
rect 20043 1503 21235 1559
rect 21291 1503 21310 1559
rect 33 1498 21310 1503
rect 4056 804 4122 807
rect 6552 804 6618 807
rect 9048 804 9114 807
rect 11544 804 11610 807
rect 14040 804 14106 807
rect 16536 804 16602 807
rect 19032 804 19098 807
rect 21528 804 21594 807
rect 0 802 21887 804
rect 0 746 4061 802
rect 4117 746 6557 802
rect 6613 746 9053 802
rect 9109 746 11549 802
rect 11605 746 14045 802
rect 14101 746 16541 802
rect 16597 746 19037 802
rect 19093 746 21533 802
rect 21589 746 21887 802
rect 0 744 21887 746
rect 4056 741 4122 744
rect 6552 741 6618 744
rect 9048 741 9114 744
rect 11544 741 11610 744
rect 14040 741 14106 744
rect 16536 741 16602 744
rect 19032 741 19098 744
rect 21528 741 21594 744
rect 3460 680 3526 683
rect 5956 680 6022 683
rect 8452 680 8518 683
rect 10948 680 11014 683
rect 13444 680 13510 683
rect 15940 680 16006 683
rect 18436 680 18502 683
rect 20932 680 20998 683
rect 0 678 21887 680
rect 0 622 3465 678
rect 3521 622 5961 678
rect 6017 622 8457 678
rect 8513 622 10953 678
rect 11009 622 13449 678
rect 13505 622 15945 678
rect 16001 622 18441 678
rect 18497 622 20937 678
rect 20993 622 21887 678
rect 0 620 21887 622
rect 3460 617 3526 620
rect 5956 617 6022 620
rect 8452 617 8518 620
rect 10948 617 11014 620
rect 13444 617 13510 620
rect 15940 617 16006 620
rect 18436 617 18502 620
rect 20932 617 20998 620
rect 2808 556 2874 559
rect 5304 556 5370 559
rect 7800 556 7866 559
rect 10296 556 10362 559
rect 12792 556 12858 559
rect 15288 556 15354 559
rect 17784 556 17850 559
rect 20280 556 20346 559
rect 0 554 21887 556
rect 0 498 2813 554
rect 2869 498 5309 554
rect 5365 498 7805 554
rect 7861 498 10301 554
rect 10357 498 12797 554
rect 12853 498 15293 554
rect 15349 498 17789 554
rect 17845 498 20285 554
rect 20341 498 21887 554
rect 0 496 21887 498
rect 2808 493 2874 496
rect 5304 493 5370 496
rect 7800 493 7866 496
rect 10296 493 10362 496
rect 12792 493 12858 496
rect 15288 493 15354 496
rect 17784 493 17850 496
rect 20280 493 20346 496
rect 2212 432 2278 435
rect 4708 432 4774 435
rect 7204 432 7270 435
rect 9700 432 9766 435
rect 12196 432 12262 435
rect 14692 432 14758 435
rect 17188 432 17254 435
rect 19684 432 19750 435
rect 0 430 21887 432
rect 0 374 2217 430
rect 2273 374 4713 430
rect 4769 374 7209 430
rect 7265 374 9705 430
rect 9761 374 12201 430
rect 12257 374 14697 430
rect 14753 374 17193 430
rect 17249 374 19689 430
rect 19745 374 21887 430
rect 0 372 21887 374
rect 2212 369 2278 372
rect 4708 369 4774 372
rect 7204 369 7270 372
rect 9700 369 9766 372
rect 12196 369 12262 372
rect 14692 369 14758 372
rect 17188 369 17254 372
rect 19684 369 19750 372
rect 1980 278 2046 281
rect 3040 278 3106 281
rect 3228 278 3294 281
rect 4288 278 4354 281
rect 1980 276 4354 278
rect 1980 220 1985 276
rect 2041 220 3045 276
rect 3101 220 3233 276
rect 3289 220 4293 276
rect 4349 220 4354 276
rect 1980 218 4354 220
rect 1980 215 2046 218
rect 3040 215 3106 218
rect 3228 215 3294 218
rect 4288 215 4354 218
rect 4476 278 4542 281
rect 5536 278 5602 281
rect 5724 278 5790 281
rect 6784 278 6850 281
rect 4476 276 6850 278
rect 4476 220 4481 276
rect 4537 220 5541 276
rect 5597 220 5729 276
rect 5785 220 6789 276
rect 6845 220 6850 276
rect 4476 218 6850 220
rect 4476 215 4542 218
rect 5536 215 5602 218
rect 5724 215 5790 218
rect 6784 215 6850 218
rect 6972 278 7038 281
rect 8032 278 8098 281
rect 8220 278 8286 281
rect 9280 278 9346 281
rect 6972 276 9346 278
rect 6972 220 6977 276
rect 7033 220 8037 276
rect 8093 220 8225 276
rect 8281 220 9285 276
rect 9341 220 9346 276
rect 6972 218 9346 220
rect 6972 215 7038 218
rect 8032 215 8098 218
rect 8220 215 8286 218
rect 9280 215 9346 218
rect 9468 278 9534 281
rect 10528 278 10594 281
rect 10716 278 10782 281
rect 11776 278 11842 281
rect 9468 276 11842 278
rect 9468 220 9473 276
rect 9529 220 10533 276
rect 10589 220 10721 276
rect 10777 220 11781 276
rect 11837 220 11842 276
rect 9468 218 11842 220
rect 9468 215 9534 218
rect 10528 215 10594 218
rect 10716 215 10782 218
rect 11776 215 11842 218
rect 11964 278 12030 281
rect 13024 278 13090 281
rect 13212 278 13278 281
rect 14272 278 14338 281
rect 11964 276 14338 278
rect 11964 220 11969 276
rect 12025 220 13029 276
rect 13085 220 13217 276
rect 13273 220 14277 276
rect 14333 220 14338 276
rect 11964 218 14338 220
rect 11964 215 12030 218
rect 13024 215 13090 218
rect 13212 215 13278 218
rect 14272 215 14338 218
rect 14460 278 14526 281
rect 15520 278 15586 281
rect 15708 278 15774 281
rect 16768 278 16834 281
rect 14460 276 16834 278
rect 14460 220 14465 276
rect 14521 220 15525 276
rect 15581 220 15713 276
rect 15769 220 16773 276
rect 16829 220 16834 276
rect 14460 218 16834 220
rect 14460 215 14526 218
rect 15520 215 15586 218
rect 15708 215 15774 218
rect 16768 215 16834 218
rect 16956 278 17022 281
rect 18016 278 18082 281
rect 18204 278 18270 281
rect 19264 278 19330 281
rect 16956 276 19330 278
rect 16956 220 16961 276
rect 17017 220 18021 276
rect 18077 220 18209 276
rect 18265 220 19269 276
rect 19325 220 19330 276
rect 16956 218 19330 220
rect 16956 215 17022 218
rect 18016 215 18082 218
rect 18204 215 18270 218
rect 19264 215 19330 218
rect 19452 278 19518 281
rect 20512 278 20578 281
rect 20700 278 20766 281
rect 21760 278 21826 281
rect 19452 276 21826 278
rect 19452 220 19457 276
rect 19513 220 20517 276
rect 20573 220 20705 276
rect 20761 220 21765 276
rect 21821 220 21826 276
rect 19452 218 21826 220
rect 19452 215 19518 218
rect 20512 215 20578 218
rect 20700 215 20766 218
rect 21760 215 21826 218
rect 2444 154 2510 157
rect 2576 154 2642 157
rect 3692 154 3758 157
rect 3824 154 3890 157
rect 2444 152 3890 154
rect 2444 96 2449 152
rect 2505 96 2581 152
rect 2637 96 3697 152
rect 3753 96 3829 152
rect 3885 96 3890 152
rect 2444 94 3890 96
rect 2444 91 2510 94
rect 2576 91 2642 94
rect 3692 91 3758 94
rect 3824 91 3890 94
rect 4940 154 5006 157
rect 5072 154 5138 157
rect 6188 154 6254 157
rect 6320 154 6386 157
rect 4940 152 6386 154
rect 4940 96 4945 152
rect 5001 96 5077 152
rect 5133 96 6193 152
rect 6249 96 6325 152
rect 6381 96 6386 152
rect 4940 94 6386 96
rect 4940 91 5006 94
rect 5072 91 5138 94
rect 6188 91 6254 94
rect 6320 91 6386 94
rect 7436 154 7502 157
rect 7568 154 7634 157
rect 8684 154 8750 157
rect 8816 154 8882 157
rect 7436 152 8882 154
rect 7436 96 7441 152
rect 7497 96 7573 152
rect 7629 96 8689 152
rect 8745 96 8821 152
rect 8877 96 8882 152
rect 7436 94 8882 96
rect 7436 91 7502 94
rect 7568 91 7634 94
rect 8684 91 8750 94
rect 8816 91 8882 94
rect 9932 154 9998 157
rect 10064 154 10130 157
rect 11180 154 11246 157
rect 11312 154 11378 157
rect 9932 152 11378 154
rect 9932 96 9937 152
rect 9993 96 10069 152
rect 10125 96 11185 152
rect 11241 96 11317 152
rect 11373 96 11378 152
rect 9932 94 11378 96
rect 9932 91 9998 94
rect 10064 91 10130 94
rect 11180 91 11246 94
rect 11312 91 11378 94
rect 12428 154 12494 157
rect 12560 154 12626 157
rect 13676 154 13742 157
rect 13808 154 13874 157
rect 12428 152 13874 154
rect 12428 96 12433 152
rect 12489 96 12565 152
rect 12621 96 13681 152
rect 13737 96 13813 152
rect 13869 96 13874 152
rect 12428 94 13874 96
rect 12428 91 12494 94
rect 12560 91 12626 94
rect 13676 91 13742 94
rect 13808 91 13874 94
rect 14924 154 14990 157
rect 15056 154 15122 157
rect 16172 154 16238 157
rect 16304 154 16370 157
rect 14924 152 16370 154
rect 14924 96 14929 152
rect 14985 96 15061 152
rect 15117 96 16177 152
rect 16233 96 16309 152
rect 16365 96 16370 152
rect 14924 94 16370 96
rect 14924 91 14990 94
rect 15056 91 15122 94
rect 16172 91 16238 94
rect 16304 91 16370 94
rect 17420 154 17486 157
rect 17552 154 17618 157
rect 18668 154 18734 157
rect 18800 154 18866 157
rect 17420 152 18866 154
rect 17420 96 17425 152
rect 17481 96 17557 152
rect 17613 96 18673 152
rect 18729 96 18805 152
rect 18861 96 18866 152
rect 17420 94 18866 96
rect 17420 91 17486 94
rect 17552 91 17618 94
rect 18668 91 18734 94
rect 18800 91 18866 94
rect 19916 154 19982 157
rect 20048 154 20114 157
rect 21164 154 21230 157
rect 21296 154 21362 157
rect 19916 152 21362 154
rect 19916 96 19921 152
rect 19977 96 20053 152
rect 20109 96 21169 152
rect 21225 96 21301 152
rect 21357 96 21362 152
rect 19916 94 21362 96
rect 19916 91 19982 94
rect 20048 91 20114 94
rect 21164 91 21230 94
rect 21296 91 21362 94
use subbyte2_column_mux_0  subbyte2_column_mux_0_0
timestamp 1543373571
transform -1 0 21887 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_1
timestamp 1543373571
transform 1 0 20639 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_2
timestamp 1543373571
transform -1 0 20639 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_3
timestamp 1543373571
transform 1 0 19391 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_4
timestamp 1543373571
transform -1 0 19391 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_5
timestamp 1543373571
transform 1 0 18143 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_6
timestamp 1543373571
transform -1 0 18143 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_7
timestamp 1543373571
transform 1 0 16895 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_8
timestamp 1543373571
transform -1 0 16895 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_9
timestamp 1543373571
transform 1 0 15647 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_10
timestamp 1543373571
transform -1 0 15647 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_11
timestamp 1543373571
transform 1 0 14399 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_12
timestamp 1543373571
transform -1 0 14399 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_13
timestamp 1543373571
transform 1 0 13151 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_14
timestamp 1543373571
transform -1 0 13151 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_15
timestamp 1543373571
transform 1 0 11903 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_16
timestamp 1543373571
transform -1 0 11903 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_17
timestamp 1543373571
transform 1 0 10655 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_18
timestamp 1543373571
transform -1 0 10655 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_19
timestamp 1543373571
transform 1 0 9407 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_20
timestamp 1543373571
transform -1 0 9407 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_21
timestamp 1543373571
transform 1 0 8159 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_22
timestamp 1543373571
transform -1 0 8159 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_23
timestamp 1543373571
transform 1 0 6911 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_24
timestamp 1543373571
transform -1 0 6911 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_25
timestamp 1543373571
transform 1 0 5663 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_26
timestamp 1543373571
transform -1 0 5663 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_27
timestamp 1543373571
transform 1 0 4415 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_28
timestamp 1543373571
transform -1 0 4415 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_29
timestamp 1543373571
transform 1 0 3167 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_30
timestamp 1543373571
transform -1 0 3167 0 1 868
box 65 0 675 1316
use subbyte2_column_mux_0  subbyte2_column_mux_0_31
timestamp 1543373571
transform 1 0 1919 0 1 868
box 65 0 675 1316
<< labels >>
rlabel metal3 s 0 372 21887 432 4 sel_0
port 3 nsew
rlabel metal3 s 0 496 21887 556 4 sel_1
port 5 nsew
rlabel metal3 s 0 620 21887 680 4 sel_2
port 7 nsew
rlabel metal3 s 0 744 21887 804 4 sel_3
port 9 nsew
rlabel metal1 s 1999 248 2027 868 4 bl_out_0
port 11 nsew
rlabel metal1 s 2463 124 2491 868 4 br_out_0
port 13 nsew
rlabel metal1 s 4495 248 4523 868 4 bl_out_1
port 15 nsew
rlabel metal1 s 4959 124 4987 868 4 br_out_1
port 17 nsew
rlabel metal1 s 6991 248 7019 868 4 bl_out_2
port 19 nsew
rlabel metal1 s 7455 124 7483 868 4 br_out_2
port 21 nsew
rlabel metal1 s 9487 248 9515 868 4 bl_out_3
port 23 nsew
rlabel metal1 s 9951 124 9979 868 4 br_out_3
port 25 nsew
rlabel metal1 s 11983 248 12011 868 4 bl_out_4
port 27 nsew
rlabel metal1 s 12447 124 12475 868 4 br_out_4
port 29 nsew
rlabel metal1 s 14479 248 14507 868 4 bl_out_5
port 31 nsew
rlabel metal1 s 14943 124 14971 868 4 br_out_5
port 33 nsew
rlabel metal1 s 16975 248 17003 868 4 bl_out_6
port 35 nsew
rlabel metal1 s 17439 124 17467 868 4 br_out_6
port 37 nsew
rlabel metal1 s 19471 248 19499 868 4 bl_out_7
port 39 nsew
rlabel metal1 s 19935 124 19963 868 4 br_out_7
port 41 nsew
rlabel metal3 s 33 1498 21310 1564 4 gnd
port 43 nsew
rlabel metal1 s 1999 2128 2027 2184 4 bl_0
port 45 nsew
rlabel metal1 s 2463 2128 2491 2184 4 br_0
port 47 nsew
rlabel metal1 s 3059 2128 3087 2184 4 bl_1
port 49 nsew
rlabel metal1 s 2595 2128 2623 2184 4 br_1
port 51 nsew
rlabel metal1 s 3247 2128 3275 2184 4 bl_2
port 53 nsew
rlabel metal1 s 3711 2128 3739 2184 4 br_2
port 55 nsew
rlabel metal1 s 4307 2128 4335 2184 4 bl_3
port 57 nsew
rlabel metal1 s 3843 2128 3871 2184 4 br_3
port 59 nsew
rlabel metal1 s 4495 2128 4523 2184 4 bl_4
port 61 nsew
rlabel metal1 s 4959 2128 4987 2184 4 br_4
port 63 nsew
rlabel metal1 s 5555 2128 5583 2184 4 bl_5
port 65 nsew
rlabel metal1 s 5091 2128 5119 2184 4 br_5
port 67 nsew
rlabel metal1 s 5743 2128 5771 2184 4 bl_6
port 69 nsew
rlabel metal1 s 6207 2128 6235 2184 4 br_6
port 71 nsew
rlabel metal1 s 6803 2128 6831 2184 4 bl_7
port 73 nsew
rlabel metal1 s 6339 2128 6367 2184 4 br_7
port 75 nsew
rlabel metal1 s 6991 2128 7019 2184 4 bl_8
port 77 nsew
rlabel metal1 s 7455 2128 7483 2184 4 br_8
port 79 nsew
rlabel metal1 s 8051 2128 8079 2184 4 bl_9
port 81 nsew
rlabel metal1 s 7587 2128 7615 2184 4 br_9
port 83 nsew
rlabel metal1 s 8239 2128 8267 2184 4 bl_10
port 85 nsew
rlabel metal1 s 8703 2128 8731 2184 4 br_10
port 87 nsew
rlabel metal1 s 9299 2128 9327 2184 4 bl_11
port 89 nsew
rlabel metal1 s 8835 2128 8863 2184 4 br_11
port 91 nsew
rlabel metal1 s 9487 2128 9515 2184 4 bl_12
port 93 nsew
rlabel metal1 s 9951 2128 9979 2184 4 br_12
port 95 nsew
rlabel metal1 s 10547 2128 10575 2184 4 bl_13
port 97 nsew
rlabel metal1 s 10083 2128 10111 2184 4 br_13
port 99 nsew
rlabel metal1 s 10735 2128 10763 2184 4 bl_14
port 101 nsew
rlabel metal1 s 11199 2128 11227 2184 4 br_14
port 103 nsew
rlabel metal1 s 11795 2128 11823 2184 4 bl_15
port 105 nsew
rlabel metal1 s 11331 2128 11359 2184 4 br_15
port 107 nsew
rlabel metal1 s 11983 2128 12011 2184 4 bl_16
port 109 nsew
rlabel metal1 s 12447 2128 12475 2184 4 br_16
port 111 nsew
rlabel metal1 s 13043 2128 13071 2184 4 bl_17
port 113 nsew
rlabel metal1 s 12579 2128 12607 2184 4 br_17
port 115 nsew
rlabel metal1 s 13231 2128 13259 2184 4 bl_18
port 117 nsew
rlabel metal1 s 13695 2128 13723 2184 4 br_18
port 119 nsew
rlabel metal1 s 14291 2128 14319 2184 4 bl_19
port 121 nsew
rlabel metal1 s 13827 2128 13855 2184 4 br_19
port 123 nsew
rlabel metal1 s 14479 2128 14507 2184 4 bl_20
port 125 nsew
rlabel metal1 s 14943 2128 14971 2184 4 br_20
port 127 nsew
rlabel metal1 s 15539 2128 15567 2184 4 bl_21
port 129 nsew
rlabel metal1 s 15075 2128 15103 2184 4 br_21
port 131 nsew
rlabel metal1 s 15727 2128 15755 2184 4 bl_22
port 133 nsew
rlabel metal1 s 16191 2128 16219 2184 4 br_22
port 135 nsew
rlabel metal1 s 16787 2128 16815 2184 4 bl_23
port 137 nsew
rlabel metal1 s 16323 2128 16351 2184 4 br_23
port 139 nsew
rlabel metal1 s 16975 2128 17003 2184 4 bl_24
port 141 nsew
rlabel metal1 s 17439 2128 17467 2184 4 br_24
port 143 nsew
rlabel metal1 s 18035 2128 18063 2184 4 bl_25
port 145 nsew
rlabel metal1 s 17571 2128 17599 2184 4 br_25
port 147 nsew
rlabel metal1 s 18223 2128 18251 2184 4 bl_26
port 149 nsew
rlabel metal1 s 18687 2128 18715 2184 4 br_26
port 151 nsew
rlabel metal1 s 19283 2128 19311 2184 4 bl_27
port 153 nsew
rlabel metal1 s 18819 2128 18847 2184 4 br_27
port 155 nsew
rlabel metal1 s 19471 2128 19499 2184 4 bl_28
port 157 nsew
rlabel metal1 s 19935 2128 19963 2184 4 br_28
port 159 nsew
rlabel metal1 s 20531 2128 20559 2184 4 bl_29
port 161 nsew
rlabel metal1 s 20067 2128 20095 2184 4 br_29
port 163 nsew
rlabel metal1 s 20719 2128 20747 2184 4 bl_30
port 165 nsew
rlabel metal1 s 21183 2128 21211 2184 4 br_30
port 167 nsew
rlabel metal1 s 21779 2128 21807 2184 4 bl_31
port 169 nsew
rlabel metal1 s 21315 2128 21343 2184 4 br_31
port 171 nsew
<< properties >>
string FIXED_BBOX 0 0 19968 87
<< end >>
