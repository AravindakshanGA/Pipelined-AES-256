magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 1988 2731
<< nwell >>
rect -36 679 728 1471
<< pwell >>
rect 28 159 554 329
rect 28 25 658 159
<< scnmos >>
rect 114 51 144 303
rect 222 51 252 303
rect 330 51 360 303
rect 438 51 468 303
<< scpmos >>
rect 114 963 144 1363
rect 222 963 252 1363
rect 330 963 360 1363
rect 438 963 468 1363
<< ndiff >>
rect 54 194 114 303
rect 54 160 62 194
rect 96 160 114 194
rect 54 51 114 160
rect 144 194 222 303
rect 144 160 166 194
rect 200 160 222 194
rect 144 51 222 160
rect 252 194 330 303
rect 252 160 274 194
rect 308 160 330 194
rect 252 51 330 160
rect 360 194 438 303
rect 360 160 382 194
rect 416 160 438 194
rect 360 51 438 160
rect 468 194 528 303
rect 468 160 486 194
rect 520 160 528 194
rect 468 51 528 160
<< pdiff >>
rect 54 1180 114 1363
rect 54 1146 62 1180
rect 96 1146 114 1180
rect 54 963 114 1146
rect 144 1180 222 1363
rect 144 1146 166 1180
rect 200 1146 222 1180
rect 144 963 222 1146
rect 252 1180 330 1363
rect 252 1146 274 1180
rect 308 1146 330 1180
rect 252 963 330 1146
rect 360 1180 438 1363
rect 360 1146 382 1180
rect 416 1146 438 1180
rect 360 963 438 1146
rect 468 1180 528 1363
rect 468 1146 486 1180
rect 520 1146 528 1180
rect 468 963 528 1146
<< ndiffc >>
rect 62 160 96 194
rect 166 160 200 194
rect 274 160 308 194
rect 382 160 416 194
rect 486 160 520 194
<< pdiffc >>
rect 62 1146 96 1180
rect 166 1146 200 1180
rect 274 1146 308 1180
rect 382 1146 416 1180
rect 486 1146 520 1180
<< psubdiff >>
rect 582 109 632 133
rect 582 75 590 109
rect 624 75 632 109
rect 582 51 632 75
<< nsubdiff >>
rect 582 1326 632 1350
rect 582 1292 590 1326
rect 624 1292 632 1326
rect 582 1268 632 1292
<< psubdiffcont >>
rect 590 75 624 109
<< nsubdiffcont >>
rect 590 1292 624 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 330 1363 360 1389
rect 438 1363 468 1389
rect 114 937 144 963
rect 222 937 252 963
rect 330 937 360 963
rect 438 937 468 963
rect 114 907 468 937
rect 114 703 144 907
rect 48 687 144 703
rect 48 653 64 687
rect 98 653 144 687
rect 48 637 144 653
rect 114 359 144 637
rect 114 329 468 359
rect 114 303 144 329
rect 222 303 252 329
rect 330 303 360 329
rect 438 303 468 329
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
<< polycont >>
rect 64 653 98 687
<< locali >>
rect 0 1397 692 1431
rect 62 1180 96 1397
rect 62 1130 96 1146
rect 166 1180 200 1196
rect 166 1096 200 1146
rect 274 1180 308 1397
rect 274 1130 308 1146
rect 382 1180 416 1196
rect 382 1096 416 1146
rect 486 1180 520 1397
rect 590 1326 624 1397
rect 590 1276 624 1292
rect 486 1130 520 1146
rect 166 1062 416 1096
rect 64 687 98 703
rect 64 637 98 653
rect 274 687 308 1062
rect 274 653 325 687
rect 274 278 308 653
rect 166 244 416 278
rect 62 194 96 210
rect 62 17 96 160
rect 166 194 200 244
rect 166 144 200 160
rect 274 194 308 210
rect 274 17 308 160
rect 382 194 416 244
rect 382 144 416 160
rect 486 194 520 210
rect 486 17 520 160
rect 590 109 624 125
rect 590 17 624 75
rect 0 -17 692 17
<< labels >>
rlabel locali s 81 670 81 670 4 A
port 1 nsew
rlabel locali s 308 670 308 670 4 Z
port 2 nsew
rlabel locali s 346 0 346 0 4 gnd
port 3 nsew
rlabel locali s 346 1414 346 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 692 1079
<< end >>
