magic
tech sky130A
magscale 1 2
timestamp 1543374230
<< checkpaint >>
rect -1260 -1260 69080 53998
<< dnwell >>
rect 1608 1608 66212 51130
<< nwell >>
rect 1524 51046 66296 51214
rect 1524 1692 1692 51046
rect 66128 1692 66296 51046
rect 1524 1524 66296 1692
<< nsubdiff >>
rect 1919 51147 1969 51171
rect 1919 51113 1927 51147
rect 1961 51113 1969 51147
rect 1919 51089 1969 51113
rect 2255 51147 2305 51171
rect 2255 51113 2263 51147
rect 2297 51113 2305 51147
rect 2255 51089 2305 51113
rect 2591 51147 2641 51171
rect 2591 51113 2599 51147
rect 2633 51113 2641 51147
rect 2591 51089 2641 51113
rect 2927 51147 2977 51171
rect 2927 51113 2935 51147
rect 2969 51113 2977 51147
rect 2927 51089 2977 51113
rect 3263 51147 3313 51171
rect 3263 51113 3271 51147
rect 3305 51113 3313 51147
rect 3263 51089 3313 51113
rect 3599 51147 3649 51171
rect 3599 51113 3607 51147
rect 3641 51113 3649 51147
rect 3599 51089 3649 51113
rect 3935 51147 3985 51171
rect 3935 51113 3943 51147
rect 3977 51113 3985 51147
rect 3935 51089 3985 51113
rect 4271 51147 4321 51171
rect 4271 51113 4279 51147
rect 4313 51113 4321 51147
rect 4271 51089 4321 51113
rect 4607 51147 4657 51171
rect 4607 51113 4615 51147
rect 4649 51113 4657 51147
rect 4607 51089 4657 51113
rect 4943 51147 4993 51171
rect 4943 51113 4951 51147
rect 4985 51113 4993 51147
rect 4943 51089 4993 51113
rect 5279 51147 5329 51171
rect 5279 51113 5287 51147
rect 5321 51113 5329 51147
rect 5279 51089 5329 51113
rect 5615 51147 5665 51171
rect 5615 51113 5623 51147
rect 5657 51113 5665 51147
rect 5615 51089 5665 51113
rect 5951 51147 6001 51171
rect 5951 51113 5959 51147
rect 5993 51113 6001 51147
rect 5951 51089 6001 51113
rect 6287 51147 6337 51171
rect 6287 51113 6295 51147
rect 6329 51113 6337 51147
rect 6287 51089 6337 51113
rect 6623 51147 6673 51171
rect 6623 51113 6631 51147
rect 6665 51113 6673 51147
rect 6623 51089 6673 51113
rect 6959 51147 7009 51171
rect 6959 51113 6967 51147
rect 7001 51113 7009 51147
rect 6959 51089 7009 51113
rect 7295 51147 7345 51171
rect 7295 51113 7303 51147
rect 7337 51113 7345 51147
rect 7295 51089 7345 51113
rect 7631 51147 7681 51171
rect 7631 51113 7639 51147
rect 7673 51113 7681 51147
rect 7631 51089 7681 51113
rect 7967 51147 8017 51171
rect 7967 51113 7975 51147
rect 8009 51113 8017 51147
rect 7967 51089 8017 51113
rect 8303 51147 8353 51171
rect 8303 51113 8311 51147
rect 8345 51113 8353 51147
rect 8303 51089 8353 51113
rect 8639 51147 8689 51171
rect 8639 51113 8647 51147
rect 8681 51113 8689 51147
rect 8639 51089 8689 51113
rect 8975 51147 9025 51171
rect 8975 51113 8983 51147
rect 9017 51113 9025 51147
rect 8975 51089 9025 51113
rect 9311 51147 9361 51171
rect 9311 51113 9319 51147
rect 9353 51113 9361 51147
rect 9311 51089 9361 51113
rect 9647 51147 9697 51171
rect 9647 51113 9655 51147
rect 9689 51113 9697 51147
rect 9647 51089 9697 51113
rect 9983 51147 10033 51171
rect 9983 51113 9991 51147
rect 10025 51113 10033 51147
rect 9983 51089 10033 51113
rect 10319 51147 10369 51171
rect 10319 51113 10327 51147
rect 10361 51113 10369 51147
rect 10319 51089 10369 51113
rect 10655 51147 10705 51171
rect 10655 51113 10663 51147
rect 10697 51113 10705 51147
rect 10655 51089 10705 51113
rect 10991 51147 11041 51171
rect 10991 51113 10999 51147
rect 11033 51113 11041 51147
rect 10991 51089 11041 51113
rect 11327 51147 11377 51171
rect 11327 51113 11335 51147
rect 11369 51113 11377 51147
rect 11327 51089 11377 51113
rect 11663 51147 11713 51171
rect 11663 51113 11671 51147
rect 11705 51113 11713 51147
rect 11663 51089 11713 51113
rect 11999 51147 12049 51171
rect 11999 51113 12007 51147
rect 12041 51113 12049 51147
rect 11999 51089 12049 51113
rect 12335 51147 12385 51171
rect 12335 51113 12343 51147
rect 12377 51113 12385 51147
rect 12335 51089 12385 51113
rect 12671 51147 12721 51171
rect 12671 51113 12679 51147
rect 12713 51113 12721 51147
rect 12671 51089 12721 51113
rect 13007 51147 13057 51171
rect 13007 51113 13015 51147
rect 13049 51113 13057 51147
rect 13007 51089 13057 51113
rect 13343 51147 13393 51171
rect 13343 51113 13351 51147
rect 13385 51113 13393 51147
rect 13343 51089 13393 51113
rect 13679 51147 13729 51171
rect 13679 51113 13687 51147
rect 13721 51113 13729 51147
rect 13679 51089 13729 51113
rect 14015 51147 14065 51171
rect 14015 51113 14023 51147
rect 14057 51113 14065 51147
rect 14015 51089 14065 51113
rect 14351 51147 14401 51171
rect 14351 51113 14359 51147
rect 14393 51113 14401 51147
rect 14351 51089 14401 51113
rect 14687 51147 14737 51171
rect 14687 51113 14695 51147
rect 14729 51113 14737 51147
rect 14687 51089 14737 51113
rect 15023 51147 15073 51171
rect 15023 51113 15031 51147
rect 15065 51113 15073 51147
rect 15023 51089 15073 51113
rect 15359 51147 15409 51171
rect 15359 51113 15367 51147
rect 15401 51113 15409 51147
rect 15359 51089 15409 51113
rect 15695 51147 15745 51171
rect 15695 51113 15703 51147
rect 15737 51113 15745 51147
rect 15695 51089 15745 51113
rect 16031 51147 16081 51171
rect 16031 51113 16039 51147
rect 16073 51113 16081 51147
rect 16031 51089 16081 51113
rect 16367 51147 16417 51171
rect 16367 51113 16375 51147
rect 16409 51113 16417 51147
rect 16367 51089 16417 51113
rect 16703 51147 16753 51171
rect 16703 51113 16711 51147
rect 16745 51113 16753 51147
rect 16703 51089 16753 51113
rect 17039 51147 17089 51171
rect 17039 51113 17047 51147
rect 17081 51113 17089 51147
rect 17039 51089 17089 51113
rect 17375 51147 17425 51171
rect 17375 51113 17383 51147
rect 17417 51113 17425 51147
rect 17375 51089 17425 51113
rect 17711 51147 17761 51171
rect 17711 51113 17719 51147
rect 17753 51113 17761 51147
rect 17711 51089 17761 51113
rect 18047 51147 18097 51171
rect 18047 51113 18055 51147
rect 18089 51113 18097 51147
rect 18047 51089 18097 51113
rect 18383 51147 18433 51171
rect 18383 51113 18391 51147
rect 18425 51113 18433 51147
rect 18383 51089 18433 51113
rect 18719 51147 18769 51171
rect 18719 51113 18727 51147
rect 18761 51113 18769 51147
rect 18719 51089 18769 51113
rect 19055 51147 19105 51171
rect 19055 51113 19063 51147
rect 19097 51113 19105 51147
rect 19055 51089 19105 51113
rect 19391 51147 19441 51171
rect 19391 51113 19399 51147
rect 19433 51113 19441 51147
rect 19391 51089 19441 51113
rect 19727 51147 19777 51171
rect 19727 51113 19735 51147
rect 19769 51113 19777 51147
rect 19727 51089 19777 51113
rect 20063 51147 20113 51171
rect 20063 51113 20071 51147
rect 20105 51113 20113 51147
rect 20063 51089 20113 51113
rect 20399 51147 20449 51171
rect 20399 51113 20407 51147
rect 20441 51113 20449 51147
rect 20399 51089 20449 51113
rect 20735 51147 20785 51171
rect 20735 51113 20743 51147
rect 20777 51113 20785 51147
rect 20735 51089 20785 51113
rect 21071 51147 21121 51171
rect 21071 51113 21079 51147
rect 21113 51113 21121 51147
rect 21071 51089 21121 51113
rect 21407 51147 21457 51171
rect 21407 51113 21415 51147
rect 21449 51113 21457 51147
rect 21407 51089 21457 51113
rect 21743 51147 21793 51171
rect 21743 51113 21751 51147
rect 21785 51113 21793 51147
rect 21743 51089 21793 51113
rect 22079 51147 22129 51171
rect 22079 51113 22087 51147
rect 22121 51113 22129 51147
rect 22079 51089 22129 51113
rect 22415 51147 22465 51171
rect 22415 51113 22423 51147
rect 22457 51113 22465 51147
rect 22415 51089 22465 51113
rect 22751 51147 22801 51171
rect 22751 51113 22759 51147
rect 22793 51113 22801 51147
rect 22751 51089 22801 51113
rect 23087 51147 23137 51171
rect 23087 51113 23095 51147
rect 23129 51113 23137 51147
rect 23087 51089 23137 51113
rect 23423 51147 23473 51171
rect 23423 51113 23431 51147
rect 23465 51113 23473 51147
rect 23423 51089 23473 51113
rect 23759 51147 23809 51171
rect 23759 51113 23767 51147
rect 23801 51113 23809 51147
rect 23759 51089 23809 51113
rect 24095 51147 24145 51171
rect 24095 51113 24103 51147
rect 24137 51113 24145 51147
rect 24095 51089 24145 51113
rect 24431 51147 24481 51171
rect 24431 51113 24439 51147
rect 24473 51113 24481 51147
rect 24431 51089 24481 51113
rect 24767 51147 24817 51171
rect 24767 51113 24775 51147
rect 24809 51113 24817 51147
rect 24767 51089 24817 51113
rect 25103 51147 25153 51171
rect 25103 51113 25111 51147
rect 25145 51113 25153 51147
rect 25103 51089 25153 51113
rect 25439 51147 25489 51171
rect 25439 51113 25447 51147
rect 25481 51113 25489 51147
rect 25439 51089 25489 51113
rect 25775 51147 25825 51171
rect 25775 51113 25783 51147
rect 25817 51113 25825 51147
rect 25775 51089 25825 51113
rect 26111 51147 26161 51171
rect 26111 51113 26119 51147
rect 26153 51113 26161 51147
rect 26111 51089 26161 51113
rect 26447 51147 26497 51171
rect 26447 51113 26455 51147
rect 26489 51113 26497 51147
rect 26447 51089 26497 51113
rect 26783 51147 26833 51171
rect 26783 51113 26791 51147
rect 26825 51113 26833 51147
rect 26783 51089 26833 51113
rect 27119 51147 27169 51171
rect 27119 51113 27127 51147
rect 27161 51113 27169 51147
rect 27119 51089 27169 51113
rect 27455 51147 27505 51171
rect 27455 51113 27463 51147
rect 27497 51113 27505 51147
rect 27455 51089 27505 51113
rect 27791 51147 27841 51171
rect 27791 51113 27799 51147
rect 27833 51113 27841 51147
rect 27791 51089 27841 51113
rect 28127 51147 28177 51171
rect 28127 51113 28135 51147
rect 28169 51113 28177 51147
rect 28127 51089 28177 51113
rect 28463 51147 28513 51171
rect 28463 51113 28471 51147
rect 28505 51113 28513 51147
rect 28463 51089 28513 51113
rect 28799 51147 28849 51171
rect 28799 51113 28807 51147
rect 28841 51113 28849 51147
rect 28799 51089 28849 51113
rect 29135 51147 29185 51171
rect 29135 51113 29143 51147
rect 29177 51113 29185 51147
rect 29135 51089 29185 51113
rect 29471 51147 29521 51171
rect 29471 51113 29479 51147
rect 29513 51113 29521 51147
rect 29471 51089 29521 51113
rect 29807 51147 29857 51171
rect 29807 51113 29815 51147
rect 29849 51113 29857 51147
rect 29807 51089 29857 51113
rect 30143 51147 30193 51171
rect 30143 51113 30151 51147
rect 30185 51113 30193 51147
rect 30143 51089 30193 51113
rect 30479 51147 30529 51171
rect 30479 51113 30487 51147
rect 30521 51113 30529 51147
rect 30479 51089 30529 51113
rect 30815 51147 30865 51171
rect 30815 51113 30823 51147
rect 30857 51113 30865 51147
rect 30815 51089 30865 51113
rect 31151 51147 31201 51171
rect 31151 51113 31159 51147
rect 31193 51113 31201 51147
rect 31151 51089 31201 51113
rect 31487 51147 31537 51171
rect 31487 51113 31495 51147
rect 31529 51113 31537 51147
rect 31487 51089 31537 51113
rect 31823 51147 31873 51171
rect 31823 51113 31831 51147
rect 31865 51113 31873 51147
rect 31823 51089 31873 51113
rect 32159 51147 32209 51171
rect 32159 51113 32167 51147
rect 32201 51113 32209 51147
rect 32159 51089 32209 51113
rect 32495 51147 32545 51171
rect 32495 51113 32503 51147
rect 32537 51113 32545 51147
rect 32495 51089 32545 51113
rect 32831 51147 32881 51171
rect 32831 51113 32839 51147
rect 32873 51113 32881 51147
rect 32831 51089 32881 51113
rect 33167 51147 33217 51171
rect 33167 51113 33175 51147
rect 33209 51113 33217 51147
rect 33167 51089 33217 51113
rect 33503 51147 33553 51171
rect 33503 51113 33511 51147
rect 33545 51113 33553 51147
rect 33503 51089 33553 51113
rect 33839 51147 33889 51171
rect 33839 51113 33847 51147
rect 33881 51113 33889 51147
rect 33839 51089 33889 51113
rect 34175 51147 34225 51171
rect 34175 51113 34183 51147
rect 34217 51113 34225 51147
rect 34175 51089 34225 51113
rect 34511 51147 34561 51171
rect 34511 51113 34519 51147
rect 34553 51113 34561 51147
rect 34511 51089 34561 51113
rect 34847 51147 34897 51171
rect 34847 51113 34855 51147
rect 34889 51113 34897 51147
rect 34847 51089 34897 51113
rect 35183 51147 35233 51171
rect 35183 51113 35191 51147
rect 35225 51113 35233 51147
rect 35183 51089 35233 51113
rect 35519 51147 35569 51171
rect 35519 51113 35527 51147
rect 35561 51113 35569 51147
rect 35519 51089 35569 51113
rect 35855 51147 35905 51171
rect 35855 51113 35863 51147
rect 35897 51113 35905 51147
rect 35855 51089 35905 51113
rect 36191 51147 36241 51171
rect 36191 51113 36199 51147
rect 36233 51113 36241 51147
rect 36191 51089 36241 51113
rect 36527 51147 36577 51171
rect 36527 51113 36535 51147
rect 36569 51113 36577 51147
rect 36527 51089 36577 51113
rect 36863 51147 36913 51171
rect 36863 51113 36871 51147
rect 36905 51113 36913 51147
rect 36863 51089 36913 51113
rect 37199 51147 37249 51171
rect 37199 51113 37207 51147
rect 37241 51113 37249 51147
rect 37199 51089 37249 51113
rect 37535 51147 37585 51171
rect 37535 51113 37543 51147
rect 37577 51113 37585 51147
rect 37535 51089 37585 51113
rect 37871 51147 37921 51171
rect 37871 51113 37879 51147
rect 37913 51113 37921 51147
rect 37871 51089 37921 51113
rect 38207 51147 38257 51171
rect 38207 51113 38215 51147
rect 38249 51113 38257 51147
rect 38207 51089 38257 51113
rect 38543 51147 38593 51171
rect 38543 51113 38551 51147
rect 38585 51113 38593 51147
rect 38543 51089 38593 51113
rect 38879 51147 38929 51171
rect 38879 51113 38887 51147
rect 38921 51113 38929 51147
rect 38879 51089 38929 51113
rect 39215 51147 39265 51171
rect 39215 51113 39223 51147
rect 39257 51113 39265 51147
rect 39215 51089 39265 51113
rect 39551 51147 39601 51171
rect 39551 51113 39559 51147
rect 39593 51113 39601 51147
rect 39551 51089 39601 51113
rect 39887 51147 39937 51171
rect 39887 51113 39895 51147
rect 39929 51113 39937 51147
rect 39887 51089 39937 51113
rect 40223 51147 40273 51171
rect 40223 51113 40231 51147
rect 40265 51113 40273 51147
rect 40223 51089 40273 51113
rect 40559 51147 40609 51171
rect 40559 51113 40567 51147
rect 40601 51113 40609 51147
rect 40559 51089 40609 51113
rect 40895 51147 40945 51171
rect 40895 51113 40903 51147
rect 40937 51113 40945 51147
rect 40895 51089 40945 51113
rect 41231 51147 41281 51171
rect 41231 51113 41239 51147
rect 41273 51113 41281 51147
rect 41231 51089 41281 51113
rect 41567 51147 41617 51171
rect 41567 51113 41575 51147
rect 41609 51113 41617 51147
rect 41567 51089 41617 51113
rect 41903 51147 41953 51171
rect 41903 51113 41911 51147
rect 41945 51113 41953 51147
rect 41903 51089 41953 51113
rect 42239 51147 42289 51171
rect 42239 51113 42247 51147
rect 42281 51113 42289 51147
rect 42239 51089 42289 51113
rect 42575 51147 42625 51171
rect 42575 51113 42583 51147
rect 42617 51113 42625 51147
rect 42575 51089 42625 51113
rect 42911 51147 42961 51171
rect 42911 51113 42919 51147
rect 42953 51113 42961 51147
rect 42911 51089 42961 51113
rect 43247 51147 43297 51171
rect 43247 51113 43255 51147
rect 43289 51113 43297 51147
rect 43247 51089 43297 51113
rect 43583 51147 43633 51171
rect 43583 51113 43591 51147
rect 43625 51113 43633 51147
rect 43583 51089 43633 51113
rect 43919 51147 43969 51171
rect 43919 51113 43927 51147
rect 43961 51113 43969 51147
rect 43919 51089 43969 51113
rect 44255 51147 44305 51171
rect 44255 51113 44263 51147
rect 44297 51113 44305 51147
rect 44255 51089 44305 51113
rect 44591 51147 44641 51171
rect 44591 51113 44599 51147
rect 44633 51113 44641 51147
rect 44591 51089 44641 51113
rect 44927 51147 44977 51171
rect 44927 51113 44935 51147
rect 44969 51113 44977 51147
rect 44927 51089 44977 51113
rect 45263 51147 45313 51171
rect 45263 51113 45271 51147
rect 45305 51113 45313 51147
rect 45263 51089 45313 51113
rect 45599 51147 45649 51171
rect 45599 51113 45607 51147
rect 45641 51113 45649 51147
rect 45599 51089 45649 51113
rect 45935 51147 45985 51171
rect 45935 51113 45943 51147
rect 45977 51113 45985 51147
rect 45935 51089 45985 51113
rect 46271 51147 46321 51171
rect 46271 51113 46279 51147
rect 46313 51113 46321 51147
rect 46271 51089 46321 51113
rect 46607 51147 46657 51171
rect 46607 51113 46615 51147
rect 46649 51113 46657 51147
rect 46607 51089 46657 51113
rect 46943 51147 46993 51171
rect 46943 51113 46951 51147
rect 46985 51113 46993 51147
rect 46943 51089 46993 51113
rect 47279 51147 47329 51171
rect 47279 51113 47287 51147
rect 47321 51113 47329 51147
rect 47279 51089 47329 51113
rect 47615 51147 47665 51171
rect 47615 51113 47623 51147
rect 47657 51113 47665 51147
rect 47615 51089 47665 51113
rect 47951 51147 48001 51171
rect 47951 51113 47959 51147
rect 47993 51113 48001 51147
rect 47951 51089 48001 51113
rect 48287 51147 48337 51171
rect 48287 51113 48295 51147
rect 48329 51113 48337 51147
rect 48287 51089 48337 51113
rect 48623 51147 48673 51171
rect 48623 51113 48631 51147
rect 48665 51113 48673 51147
rect 48623 51089 48673 51113
rect 48959 51147 49009 51171
rect 48959 51113 48967 51147
rect 49001 51113 49009 51147
rect 48959 51089 49009 51113
rect 49295 51147 49345 51171
rect 49295 51113 49303 51147
rect 49337 51113 49345 51147
rect 49295 51089 49345 51113
rect 49631 51147 49681 51171
rect 49631 51113 49639 51147
rect 49673 51113 49681 51147
rect 49631 51089 49681 51113
rect 49967 51147 50017 51171
rect 49967 51113 49975 51147
rect 50009 51113 50017 51147
rect 49967 51089 50017 51113
rect 50303 51147 50353 51171
rect 50303 51113 50311 51147
rect 50345 51113 50353 51147
rect 50303 51089 50353 51113
rect 50639 51147 50689 51171
rect 50639 51113 50647 51147
rect 50681 51113 50689 51147
rect 50639 51089 50689 51113
rect 50975 51147 51025 51171
rect 50975 51113 50983 51147
rect 51017 51113 51025 51147
rect 50975 51089 51025 51113
rect 51311 51147 51361 51171
rect 51311 51113 51319 51147
rect 51353 51113 51361 51147
rect 51311 51089 51361 51113
rect 51647 51147 51697 51171
rect 51647 51113 51655 51147
rect 51689 51113 51697 51147
rect 51647 51089 51697 51113
rect 51983 51147 52033 51171
rect 51983 51113 51991 51147
rect 52025 51113 52033 51147
rect 51983 51089 52033 51113
rect 52319 51147 52369 51171
rect 52319 51113 52327 51147
rect 52361 51113 52369 51147
rect 52319 51089 52369 51113
rect 52655 51147 52705 51171
rect 52655 51113 52663 51147
rect 52697 51113 52705 51147
rect 52655 51089 52705 51113
rect 52991 51147 53041 51171
rect 52991 51113 52999 51147
rect 53033 51113 53041 51147
rect 52991 51089 53041 51113
rect 53327 51147 53377 51171
rect 53327 51113 53335 51147
rect 53369 51113 53377 51147
rect 53327 51089 53377 51113
rect 53663 51147 53713 51171
rect 53663 51113 53671 51147
rect 53705 51113 53713 51147
rect 53663 51089 53713 51113
rect 53999 51147 54049 51171
rect 53999 51113 54007 51147
rect 54041 51113 54049 51147
rect 53999 51089 54049 51113
rect 54335 51147 54385 51171
rect 54335 51113 54343 51147
rect 54377 51113 54385 51147
rect 54335 51089 54385 51113
rect 54671 51147 54721 51171
rect 54671 51113 54679 51147
rect 54713 51113 54721 51147
rect 54671 51089 54721 51113
rect 55007 51147 55057 51171
rect 55007 51113 55015 51147
rect 55049 51113 55057 51147
rect 55007 51089 55057 51113
rect 55343 51147 55393 51171
rect 55343 51113 55351 51147
rect 55385 51113 55393 51147
rect 55343 51089 55393 51113
rect 55679 51147 55729 51171
rect 55679 51113 55687 51147
rect 55721 51113 55729 51147
rect 55679 51089 55729 51113
rect 56015 51147 56065 51171
rect 56015 51113 56023 51147
rect 56057 51113 56065 51147
rect 56015 51089 56065 51113
rect 56351 51147 56401 51171
rect 56351 51113 56359 51147
rect 56393 51113 56401 51147
rect 56351 51089 56401 51113
rect 56687 51147 56737 51171
rect 56687 51113 56695 51147
rect 56729 51113 56737 51147
rect 56687 51089 56737 51113
rect 57023 51147 57073 51171
rect 57023 51113 57031 51147
rect 57065 51113 57073 51147
rect 57023 51089 57073 51113
rect 57359 51147 57409 51171
rect 57359 51113 57367 51147
rect 57401 51113 57409 51147
rect 57359 51089 57409 51113
rect 57695 51147 57745 51171
rect 57695 51113 57703 51147
rect 57737 51113 57745 51147
rect 57695 51089 57745 51113
rect 58031 51147 58081 51171
rect 58031 51113 58039 51147
rect 58073 51113 58081 51147
rect 58031 51089 58081 51113
rect 58367 51147 58417 51171
rect 58367 51113 58375 51147
rect 58409 51113 58417 51147
rect 58367 51089 58417 51113
rect 58703 51147 58753 51171
rect 58703 51113 58711 51147
rect 58745 51113 58753 51147
rect 58703 51089 58753 51113
rect 59039 51147 59089 51171
rect 59039 51113 59047 51147
rect 59081 51113 59089 51147
rect 59039 51089 59089 51113
rect 59375 51147 59425 51171
rect 59375 51113 59383 51147
rect 59417 51113 59425 51147
rect 59375 51089 59425 51113
rect 59711 51147 59761 51171
rect 59711 51113 59719 51147
rect 59753 51113 59761 51147
rect 59711 51089 59761 51113
rect 60047 51147 60097 51171
rect 60047 51113 60055 51147
rect 60089 51113 60097 51147
rect 60047 51089 60097 51113
rect 60383 51147 60433 51171
rect 60383 51113 60391 51147
rect 60425 51113 60433 51147
rect 60383 51089 60433 51113
rect 60719 51147 60769 51171
rect 60719 51113 60727 51147
rect 60761 51113 60769 51147
rect 60719 51089 60769 51113
rect 61055 51147 61105 51171
rect 61055 51113 61063 51147
rect 61097 51113 61105 51147
rect 61055 51089 61105 51113
rect 61391 51147 61441 51171
rect 61391 51113 61399 51147
rect 61433 51113 61441 51147
rect 61391 51089 61441 51113
rect 61727 51147 61777 51171
rect 61727 51113 61735 51147
rect 61769 51113 61777 51147
rect 61727 51089 61777 51113
rect 62063 51147 62113 51171
rect 62063 51113 62071 51147
rect 62105 51113 62113 51147
rect 62063 51089 62113 51113
rect 62399 51147 62449 51171
rect 62399 51113 62407 51147
rect 62441 51113 62449 51147
rect 62399 51089 62449 51113
rect 62735 51147 62785 51171
rect 62735 51113 62743 51147
rect 62777 51113 62785 51147
rect 62735 51089 62785 51113
rect 63071 51147 63121 51171
rect 63071 51113 63079 51147
rect 63113 51113 63121 51147
rect 63071 51089 63121 51113
rect 63407 51147 63457 51171
rect 63407 51113 63415 51147
rect 63449 51113 63457 51147
rect 63407 51089 63457 51113
rect 63743 51147 63793 51171
rect 63743 51113 63751 51147
rect 63785 51113 63793 51147
rect 63743 51089 63793 51113
rect 64079 51147 64129 51171
rect 64079 51113 64087 51147
rect 64121 51113 64129 51147
rect 64079 51089 64129 51113
rect 64415 51147 64465 51171
rect 64415 51113 64423 51147
rect 64457 51113 64465 51147
rect 64415 51089 64465 51113
rect 64751 51147 64801 51171
rect 64751 51113 64759 51147
rect 64793 51113 64801 51147
rect 64751 51089 64801 51113
rect 65087 51147 65137 51171
rect 65087 51113 65095 51147
rect 65129 51113 65137 51147
rect 65087 51089 65137 51113
rect 65423 51147 65473 51171
rect 65423 51113 65431 51147
rect 65465 51113 65473 51147
rect 65423 51089 65473 51113
rect 65759 51147 65809 51171
rect 65759 51113 65767 51147
rect 65801 51113 65809 51147
rect 65759 51089 65809 51113
rect 1583 50681 1633 50705
rect 1583 50647 1591 50681
rect 1625 50647 1633 50681
rect 1583 50623 1633 50647
rect 66187 50681 66237 50705
rect 66187 50647 66195 50681
rect 66229 50647 66237 50681
rect 66187 50623 66237 50647
rect 1583 50345 1633 50369
rect 1583 50311 1591 50345
rect 1625 50311 1633 50345
rect 1583 50287 1633 50311
rect 66187 50345 66237 50369
rect 66187 50311 66195 50345
rect 66229 50311 66237 50345
rect 66187 50287 66237 50311
rect 1583 50009 1633 50033
rect 1583 49975 1591 50009
rect 1625 49975 1633 50009
rect 1583 49951 1633 49975
rect 66187 50009 66237 50033
rect 66187 49975 66195 50009
rect 66229 49975 66237 50009
rect 66187 49951 66237 49975
rect 1583 49673 1633 49697
rect 1583 49639 1591 49673
rect 1625 49639 1633 49673
rect 1583 49615 1633 49639
rect 66187 49673 66237 49697
rect 66187 49639 66195 49673
rect 66229 49639 66237 49673
rect 66187 49615 66237 49639
rect 1583 49337 1633 49361
rect 1583 49303 1591 49337
rect 1625 49303 1633 49337
rect 1583 49279 1633 49303
rect 66187 49337 66237 49361
rect 66187 49303 66195 49337
rect 66229 49303 66237 49337
rect 66187 49279 66237 49303
rect 1583 49001 1633 49025
rect 1583 48967 1591 49001
rect 1625 48967 1633 49001
rect 1583 48943 1633 48967
rect 66187 49001 66237 49025
rect 66187 48967 66195 49001
rect 66229 48967 66237 49001
rect 66187 48943 66237 48967
rect 1583 48665 1633 48689
rect 1583 48631 1591 48665
rect 1625 48631 1633 48665
rect 1583 48607 1633 48631
rect 66187 48665 66237 48689
rect 66187 48631 66195 48665
rect 66229 48631 66237 48665
rect 66187 48607 66237 48631
rect 1583 48329 1633 48353
rect 1583 48295 1591 48329
rect 1625 48295 1633 48329
rect 1583 48271 1633 48295
rect 66187 48329 66237 48353
rect 66187 48295 66195 48329
rect 66229 48295 66237 48329
rect 66187 48271 66237 48295
rect 1583 47993 1633 48017
rect 1583 47959 1591 47993
rect 1625 47959 1633 47993
rect 1583 47935 1633 47959
rect 66187 47993 66237 48017
rect 66187 47959 66195 47993
rect 66229 47959 66237 47993
rect 66187 47935 66237 47959
rect 1583 47657 1633 47681
rect 1583 47623 1591 47657
rect 1625 47623 1633 47657
rect 1583 47599 1633 47623
rect 66187 47657 66237 47681
rect 66187 47623 66195 47657
rect 66229 47623 66237 47657
rect 66187 47599 66237 47623
rect 1583 47321 1633 47345
rect 1583 47287 1591 47321
rect 1625 47287 1633 47321
rect 1583 47263 1633 47287
rect 66187 47321 66237 47345
rect 66187 47287 66195 47321
rect 66229 47287 66237 47321
rect 66187 47263 66237 47287
rect 1583 46985 1633 47009
rect 1583 46951 1591 46985
rect 1625 46951 1633 46985
rect 1583 46927 1633 46951
rect 66187 46985 66237 47009
rect 66187 46951 66195 46985
rect 66229 46951 66237 46985
rect 66187 46927 66237 46951
rect 1583 46649 1633 46673
rect 1583 46615 1591 46649
rect 1625 46615 1633 46649
rect 1583 46591 1633 46615
rect 66187 46649 66237 46673
rect 66187 46615 66195 46649
rect 66229 46615 66237 46649
rect 66187 46591 66237 46615
rect 1583 46313 1633 46337
rect 1583 46279 1591 46313
rect 1625 46279 1633 46313
rect 1583 46255 1633 46279
rect 66187 46313 66237 46337
rect 66187 46279 66195 46313
rect 66229 46279 66237 46313
rect 66187 46255 66237 46279
rect 1583 45977 1633 46001
rect 1583 45943 1591 45977
rect 1625 45943 1633 45977
rect 1583 45919 1633 45943
rect 66187 45977 66237 46001
rect 66187 45943 66195 45977
rect 66229 45943 66237 45977
rect 66187 45919 66237 45943
rect 1583 45641 1633 45665
rect 1583 45607 1591 45641
rect 1625 45607 1633 45641
rect 1583 45583 1633 45607
rect 66187 45641 66237 45665
rect 66187 45607 66195 45641
rect 66229 45607 66237 45641
rect 66187 45583 66237 45607
rect 1583 45305 1633 45329
rect 1583 45271 1591 45305
rect 1625 45271 1633 45305
rect 1583 45247 1633 45271
rect 66187 45305 66237 45329
rect 66187 45271 66195 45305
rect 66229 45271 66237 45305
rect 66187 45247 66237 45271
rect 1583 44969 1633 44993
rect 1583 44935 1591 44969
rect 1625 44935 1633 44969
rect 1583 44911 1633 44935
rect 66187 44969 66237 44993
rect 66187 44935 66195 44969
rect 66229 44935 66237 44969
rect 66187 44911 66237 44935
rect 1583 44633 1633 44657
rect 1583 44599 1591 44633
rect 1625 44599 1633 44633
rect 1583 44575 1633 44599
rect 66187 44633 66237 44657
rect 66187 44599 66195 44633
rect 66229 44599 66237 44633
rect 66187 44575 66237 44599
rect 1583 44297 1633 44321
rect 1583 44263 1591 44297
rect 1625 44263 1633 44297
rect 1583 44239 1633 44263
rect 66187 44297 66237 44321
rect 66187 44263 66195 44297
rect 66229 44263 66237 44297
rect 66187 44239 66237 44263
rect 1583 43961 1633 43985
rect 1583 43927 1591 43961
rect 1625 43927 1633 43961
rect 1583 43903 1633 43927
rect 66187 43961 66237 43985
rect 66187 43927 66195 43961
rect 66229 43927 66237 43961
rect 66187 43903 66237 43927
rect 1583 43625 1633 43649
rect 1583 43591 1591 43625
rect 1625 43591 1633 43625
rect 1583 43567 1633 43591
rect 66187 43625 66237 43649
rect 66187 43591 66195 43625
rect 66229 43591 66237 43625
rect 66187 43567 66237 43591
rect 1583 43289 1633 43313
rect 1583 43255 1591 43289
rect 1625 43255 1633 43289
rect 1583 43231 1633 43255
rect 66187 43289 66237 43313
rect 66187 43255 66195 43289
rect 66229 43255 66237 43289
rect 66187 43231 66237 43255
rect 1583 42953 1633 42977
rect 1583 42919 1591 42953
rect 1625 42919 1633 42953
rect 1583 42895 1633 42919
rect 66187 42953 66237 42977
rect 66187 42919 66195 42953
rect 66229 42919 66237 42953
rect 66187 42895 66237 42919
rect 1583 42617 1633 42641
rect 1583 42583 1591 42617
rect 1625 42583 1633 42617
rect 1583 42559 1633 42583
rect 66187 42617 66237 42641
rect 66187 42583 66195 42617
rect 66229 42583 66237 42617
rect 66187 42559 66237 42583
rect 1583 42281 1633 42305
rect 1583 42247 1591 42281
rect 1625 42247 1633 42281
rect 1583 42223 1633 42247
rect 66187 42281 66237 42305
rect 66187 42247 66195 42281
rect 66229 42247 66237 42281
rect 66187 42223 66237 42247
rect 1583 41945 1633 41969
rect 1583 41911 1591 41945
rect 1625 41911 1633 41945
rect 1583 41887 1633 41911
rect 66187 41945 66237 41969
rect 66187 41911 66195 41945
rect 66229 41911 66237 41945
rect 66187 41887 66237 41911
rect 1583 41609 1633 41633
rect 1583 41575 1591 41609
rect 1625 41575 1633 41609
rect 1583 41551 1633 41575
rect 66187 41609 66237 41633
rect 66187 41575 66195 41609
rect 66229 41575 66237 41609
rect 66187 41551 66237 41575
rect 1583 41273 1633 41297
rect 1583 41239 1591 41273
rect 1625 41239 1633 41273
rect 1583 41215 1633 41239
rect 66187 41273 66237 41297
rect 66187 41239 66195 41273
rect 66229 41239 66237 41273
rect 66187 41215 66237 41239
rect 1583 40937 1633 40961
rect 1583 40903 1591 40937
rect 1625 40903 1633 40937
rect 1583 40879 1633 40903
rect 66187 40937 66237 40961
rect 66187 40903 66195 40937
rect 66229 40903 66237 40937
rect 66187 40879 66237 40903
rect 1583 40601 1633 40625
rect 1583 40567 1591 40601
rect 1625 40567 1633 40601
rect 1583 40543 1633 40567
rect 66187 40601 66237 40625
rect 66187 40567 66195 40601
rect 66229 40567 66237 40601
rect 66187 40543 66237 40567
rect 1583 40265 1633 40289
rect 1583 40231 1591 40265
rect 1625 40231 1633 40265
rect 1583 40207 1633 40231
rect 66187 40265 66237 40289
rect 66187 40231 66195 40265
rect 66229 40231 66237 40265
rect 66187 40207 66237 40231
rect 1583 39929 1633 39953
rect 1583 39895 1591 39929
rect 1625 39895 1633 39929
rect 1583 39871 1633 39895
rect 66187 39929 66237 39953
rect 66187 39895 66195 39929
rect 66229 39895 66237 39929
rect 66187 39871 66237 39895
rect 1583 39593 1633 39617
rect 1583 39559 1591 39593
rect 1625 39559 1633 39593
rect 1583 39535 1633 39559
rect 66187 39593 66237 39617
rect 66187 39559 66195 39593
rect 66229 39559 66237 39593
rect 66187 39535 66237 39559
rect 1583 39257 1633 39281
rect 1583 39223 1591 39257
rect 1625 39223 1633 39257
rect 1583 39199 1633 39223
rect 66187 39257 66237 39281
rect 66187 39223 66195 39257
rect 66229 39223 66237 39257
rect 66187 39199 66237 39223
rect 1583 38921 1633 38945
rect 1583 38887 1591 38921
rect 1625 38887 1633 38921
rect 1583 38863 1633 38887
rect 66187 38921 66237 38945
rect 66187 38887 66195 38921
rect 66229 38887 66237 38921
rect 66187 38863 66237 38887
rect 1583 38585 1633 38609
rect 1583 38551 1591 38585
rect 1625 38551 1633 38585
rect 1583 38527 1633 38551
rect 66187 38585 66237 38609
rect 66187 38551 66195 38585
rect 66229 38551 66237 38585
rect 66187 38527 66237 38551
rect 1583 38249 1633 38273
rect 1583 38215 1591 38249
rect 1625 38215 1633 38249
rect 1583 38191 1633 38215
rect 66187 38249 66237 38273
rect 66187 38215 66195 38249
rect 66229 38215 66237 38249
rect 66187 38191 66237 38215
rect 1583 37913 1633 37937
rect 1583 37879 1591 37913
rect 1625 37879 1633 37913
rect 1583 37855 1633 37879
rect 66187 37913 66237 37937
rect 66187 37879 66195 37913
rect 66229 37879 66237 37913
rect 66187 37855 66237 37879
rect 1583 37577 1633 37601
rect 1583 37543 1591 37577
rect 1625 37543 1633 37577
rect 1583 37519 1633 37543
rect 66187 37577 66237 37601
rect 66187 37543 66195 37577
rect 66229 37543 66237 37577
rect 66187 37519 66237 37543
rect 1583 37241 1633 37265
rect 1583 37207 1591 37241
rect 1625 37207 1633 37241
rect 1583 37183 1633 37207
rect 66187 37241 66237 37265
rect 66187 37207 66195 37241
rect 66229 37207 66237 37241
rect 66187 37183 66237 37207
rect 1583 36905 1633 36929
rect 1583 36871 1591 36905
rect 1625 36871 1633 36905
rect 1583 36847 1633 36871
rect 66187 36905 66237 36929
rect 66187 36871 66195 36905
rect 66229 36871 66237 36905
rect 66187 36847 66237 36871
rect 1583 36569 1633 36593
rect 1583 36535 1591 36569
rect 1625 36535 1633 36569
rect 1583 36511 1633 36535
rect 66187 36569 66237 36593
rect 66187 36535 66195 36569
rect 66229 36535 66237 36569
rect 66187 36511 66237 36535
rect 1583 36233 1633 36257
rect 1583 36199 1591 36233
rect 1625 36199 1633 36233
rect 1583 36175 1633 36199
rect 66187 36233 66237 36257
rect 66187 36199 66195 36233
rect 66229 36199 66237 36233
rect 66187 36175 66237 36199
rect 1583 35897 1633 35921
rect 1583 35863 1591 35897
rect 1625 35863 1633 35897
rect 1583 35839 1633 35863
rect 66187 35897 66237 35921
rect 66187 35863 66195 35897
rect 66229 35863 66237 35897
rect 66187 35839 66237 35863
rect 1583 35561 1633 35585
rect 1583 35527 1591 35561
rect 1625 35527 1633 35561
rect 1583 35503 1633 35527
rect 66187 35561 66237 35585
rect 66187 35527 66195 35561
rect 66229 35527 66237 35561
rect 66187 35503 66237 35527
rect 1583 35225 1633 35249
rect 1583 35191 1591 35225
rect 1625 35191 1633 35225
rect 1583 35167 1633 35191
rect 66187 35225 66237 35249
rect 66187 35191 66195 35225
rect 66229 35191 66237 35225
rect 66187 35167 66237 35191
rect 1583 34889 1633 34913
rect 1583 34855 1591 34889
rect 1625 34855 1633 34889
rect 1583 34831 1633 34855
rect 66187 34889 66237 34913
rect 66187 34855 66195 34889
rect 66229 34855 66237 34889
rect 66187 34831 66237 34855
rect 1583 34553 1633 34577
rect 1583 34519 1591 34553
rect 1625 34519 1633 34553
rect 1583 34495 1633 34519
rect 66187 34553 66237 34577
rect 66187 34519 66195 34553
rect 66229 34519 66237 34553
rect 66187 34495 66237 34519
rect 1583 34217 1633 34241
rect 1583 34183 1591 34217
rect 1625 34183 1633 34217
rect 1583 34159 1633 34183
rect 66187 34217 66237 34241
rect 66187 34183 66195 34217
rect 66229 34183 66237 34217
rect 66187 34159 66237 34183
rect 1583 33881 1633 33905
rect 1583 33847 1591 33881
rect 1625 33847 1633 33881
rect 1583 33823 1633 33847
rect 66187 33881 66237 33905
rect 66187 33847 66195 33881
rect 66229 33847 66237 33881
rect 66187 33823 66237 33847
rect 1583 33545 1633 33569
rect 1583 33511 1591 33545
rect 1625 33511 1633 33545
rect 1583 33487 1633 33511
rect 66187 33545 66237 33569
rect 66187 33511 66195 33545
rect 66229 33511 66237 33545
rect 66187 33487 66237 33511
rect 1583 33209 1633 33233
rect 1583 33175 1591 33209
rect 1625 33175 1633 33209
rect 1583 33151 1633 33175
rect 66187 33209 66237 33233
rect 66187 33175 66195 33209
rect 66229 33175 66237 33209
rect 66187 33151 66237 33175
rect 1583 32873 1633 32897
rect 1583 32839 1591 32873
rect 1625 32839 1633 32873
rect 1583 32815 1633 32839
rect 66187 32873 66237 32897
rect 66187 32839 66195 32873
rect 66229 32839 66237 32873
rect 66187 32815 66237 32839
rect 1583 32537 1633 32561
rect 1583 32503 1591 32537
rect 1625 32503 1633 32537
rect 1583 32479 1633 32503
rect 66187 32537 66237 32561
rect 66187 32503 66195 32537
rect 66229 32503 66237 32537
rect 66187 32479 66237 32503
rect 1583 32201 1633 32225
rect 1583 32167 1591 32201
rect 1625 32167 1633 32201
rect 1583 32143 1633 32167
rect 66187 32201 66237 32225
rect 66187 32167 66195 32201
rect 66229 32167 66237 32201
rect 66187 32143 66237 32167
rect 1583 31865 1633 31889
rect 1583 31831 1591 31865
rect 1625 31831 1633 31865
rect 1583 31807 1633 31831
rect 66187 31865 66237 31889
rect 66187 31831 66195 31865
rect 66229 31831 66237 31865
rect 66187 31807 66237 31831
rect 1583 31529 1633 31553
rect 1583 31495 1591 31529
rect 1625 31495 1633 31529
rect 1583 31471 1633 31495
rect 66187 31529 66237 31553
rect 66187 31495 66195 31529
rect 66229 31495 66237 31529
rect 66187 31471 66237 31495
rect 1583 31193 1633 31217
rect 1583 31159 1591 31193
rect 1625 31159 1633 31193
rect 1583 31135 1633 31159
rect 66187 31193 66237 31217
rect 66187 31159 66195 31193
rect 66229 31159 66237 31193
rect 66187 31135 66237 31159
rect 1583 30857 1633 30881
rect 1583 30823 1591 30857
rect 1625 30823 1633 30857
rect 1583 30799 1633 30823
rect 66187 30857 66237 30881
rect 66187 30823 66195 30857
rect 66229 30823 66237 30857
rect 66187 30799 66237 30823
rect 1583 30521 1633 30545
rect 1583 30487 1591 30521
rect 1625 30487 1633 30521
rect 1583 30463 1633 30487
rect 66187 30521 66237 30545
rect 66187 30487 66195 30521
rect 66229 30487 66237 30521
rect 66187 30463 66237 30487
rect 1583 30185 1633 30209
rect 1583 30151 1591 30185
rect 1625 30151 1633 30185
rect 1583 30127 1633 30151
rect 66187 30185 66237 30209
rect 66187 30151 66195 30185
rect 66229 30151 66237 30185
rect 66187 30127 66237 30151
rect 1583 29849 1633 29873
rect 1583 29815 1591 29849
rect 1625 29815 1633 29849
rect 1583 29791 1633 29815
rect 66187 29849 66237 29873
rect 66187 29815 66195 29849
rect 66229 29815 66237 29849
rect 66187 29791 66237 29815
rect 1583 29513 1633 29537
rect 1583 29479 1591 29513
rect 1625 29479 1633 29513
rect 1583 29455 1633 29479
rect 66187 29513 66237 29537
rect 66187 29479 66195 29513
rect 66229 29479 66237 29513
rect 66187 29455 66237 29479
rect 1583 29177 1633 29201
rect 1583 29143 1591 29177
rect 1625 29143 1633 29177
rect 1583 29119 1633 29143
rect 66187 29177 66237 29201
rect 66187 29143 66195 29177
rect 66229 29143 66237 29177
rect 66187 29119 66237 29143
rect 1583 28841 1633 28865
rect 1583 28807 1591 28841
rect 1625 28807 1633 28841
rect 1583 28783 1633 28807
rect 66187 28841 66237 28865
rect 66187 28807 66195 28841
rect 66229 28807 66237 28841
rect 66187 28783 66237 28807
rect 1583 28505 1633 28529
rect 1583 28471 1591 28505
rect 1625 28471 1633 28505
rect 1583 28447 1633 28471
rect 66187 28505 66237 28529
rect 66187 28471 66195 28505
rect 66229 28471 66237 28505
rect 66187 28447 66237 28471
rect 1583 28169 1633 28193
rect 1583 28135 1591 28169
rect 1625 28135 1633 28169
rect 1583 28111 1633 28135
rect 66187 28169 66237 28193
rect 66187 28135 66195 28169
rect 66229 28135 66237 28169
rect 66187 28111 66237 28135
rect 1583 27833 1633 27857
rect 1583 27799 1591 27833
rect 1625 27799 1633 27833
rect 1583 27775 1633 27799
rect 66187 27833 66237 27857
rect 66187 27799 66195 27833
rect 66229 27799 66237 27833
rect 66187 27775 66237 27799
rect 1583 27497 1633 27521
rect 1583 27463 1591 27497
rect 1625 27463 1633 27497
rect 1583 27439 1633 27463
rect 66187 27497 66237 27521
rect 66187 27463 66195 27497
rect 66229 27463 66237 27497
rect 66187 27439 66237 27463
rect 1583 27161 1633 27185
rect 1583 27127 1591 27161
rect 1625 27127 1633 27161
rect 1583 27103 1633 27127
rect 66187 27161 66237 27185
rect 66187 27127 66195 27161
rect 66229 27127 66237 27161
rect 66187 27103 66237 27127
rect 1583 26825 1633 26849
rect 1583 26791 1591 26825
rect 1625 26791 1633 26825
rect 1583 26767 1633 26791
rect 66187 26825 66237 26849
rect 66187 26791 66195 26825
rect 66229 26791 66237 26825
rect 66187 26767 66237 26791
rect 1583 26489 1633 26513
rect 1583 26455 1591 26489
rect 1625 26455 1633 26489
rect 1583 26431 1633 26455
rect 66187 26489 66237 26513
rect 66187 26455 66195 26489
rect 66229 26455 66237 26489
rect 66187 26431 66237 26455
rect 1583 26153 1633 26177
rect 1583 26119 1591 26153
rect 1625 26119 1633 26153
rect 1583 26095 1633 26119
rect 66187 26153 66237 26177
rect 66187 26119 66195 26153
rect 66229 26119 66237 26153
rect 66187 26095 66237 26119
rect 1583 25817 1633 25841
rect 1583 25783 1591 25817
rect 1625 25783 1633 25817
rect 1583 25759 1633 25783
rect 66187 25817 66237 25841
rect 66187 25783 66195 25817
rect 66229 25783 66237 25817
rect 66187 25759 66237 25783
rect 1583 25481 1633 25505
rect 1583 25447 1591 25481
rect 1625 25447 1633 25481
rect 1583 25423 1633 25447
rect 66187 25481 66237 25505
rect 66187 25447 66195 25481
rect 66229 25447 66237 25481
rect 66187 25423 66237 25447
rect 1583 25145 1633 25169
rect 1583 25111 1591 25145
rect 1625 25111 1633 25145
rect 1583 25087 1633 25111
rect 66187 25145 66237 25169
rect 66187 25111 66195 25145
rect 66229 25111 66237 25145
rect 66187 25087 66237 25111
rect 1583 24809 1633 24833
rect 1583 24775 1591 24809
rect 1625 24775 1633 24809
rect 1583 24751 1633 24775
rect 66187 24809 66237 24833
rect 66187 24775 66195 24809
rect 66229 24775 66237 24809
rect 66187 24751 66237 24775
rect 1583 24473 1633 24497
rect 1583 24439 1591 24473
rect 1625 24439 1633 24473
rect 1583 24415 1633 24439
rect 66187 24473 66237 24497
rect 66187 24439 66195 24473
rect 66229 24439 66237 24473
rect 66187 24415 66237 24439
rect 1583 24137 1633 24161
rect 1583 24103 1591 24137
rect 1625 24103 1633 24137
rect 1583 24079 1633 24103
rect 66187 24137 66237 24161
rect 66187 24103 66195 24137
rect 66229 24103 66237 24137
rect 66187 24079 66237 24103
rect 1583 23801 1633 23825
rect 1583 23767 1591 23801
rect 1625 23767 1633 23801
rect 1583 23743 1633 23767
rect 66187 23801 66237 23825
rect 66187 23767 66195 23801
rect 66229 23767 66237 23801
rect 66187 23743 66237 23767
rect 1583 23465 1633 23489
rect 1583 23431 1591 23465
rect 1625 23431 1633 23465
rect 1583 23407 1633 23431
rect 66187 23465 66237 23489
rect 66187 23431 66195 23465
rect 66229 23431 66237 23465
rect 66187 23407 66237 23431
rect 1583 23129 1633 23153
rect 1583 23095 1591 23129
rect 1625 23095 1633 23129
rect 1583 23071 1633 23095
rect 66187 23129 66237 23153
rect 66187 23095 66195 23129
rect 66229 23095 66237 23129
rect 66187 23071 66237 23095
rect 1583 22793 1633 22817
rect 1583 22759 1591 22793
rect 1625 22759 1633 22793
rect 1583 22735 1633 22759
rect 66187 22793 66237 22817
rect 66187 22759 66195 22793
rect 66229 22759 66237 22793
rect 66187 22735 66237 22759
rect 1583 22457 1633 22481
rect 1583 22423 1591 22457
rect 1625 22423 1633 22457
rect 1583 22399 1633 22423
rect 66187 22457 66237 22481
rect 66187 22423 66195 22457
rect 66229 22423 66237 22457
rect 66187 22399 66237 22423
rect 1583 22121 1633 22145
rect 1583 22087 1591 22121
rect 1625 22087 1633 22121
rect 1583 22063 1633 22087
rect 66187 22121 66237 22145
rect 66187 22087 66195 22121
rect 66229 22087 66237 22121
rect 66187 22063 66237 22087
rect 1583 21785 1633 21809
rect 1583 21751 1591 21785
rect 1625 21751 1633 21785
rect 1583 21727 1633 21751
rect 66187 21785 66237 21809
rect 66187 21751 66195 21785
rect 66229 21751 66237 21785
rect 66187 21727 66237 21751
rect 1583 21449 1633 21473
rect 1583 21415 1591 21449
rect 1625 21415 1633 21449
rect 1583 21391 1633 21415
rect 66187 21449 66237 21473
rect 66187 21415 66195 21449
rect 66229 21415 66237 21449
rect 66187 21391 66237 21415
rect 1583 21113 1633 21137
rect 1583 21079 1591 21113
rect 1625 21079 1633 21113
rect 1583 21055 1633 21079
rect 66187 21113 66237 21137
rect 66187 21079 66195 21113
rect 66229 21079 66237 21113
rect 66187 21055 66237 21079
rect 1583 20777 1633 20801
rect 1583 20743 1591 20777
rect 1625 20743 1633 20777
rect 1583 20719 1633 20743
rect 66187 20777 66237 20801
rect 66187 20743 66195 20777
rect 66229 20743 66237 20777
rect 66187 20719 66237 20743
rect 1583 20441 1633 20465
rect 1583 20407 1591 20441
rect 1625 20407 1633 20441
rect 1583 20383 1633 20407
rect 66187 20441 66237 20465
rect 66187 20407 66195 20441
rect 66229 20407 66237 20441
rect 66187 20383 66237 20407
rect 1583 20105 1633 20129
rect 1583 20071 1591 20105
rect 1625 20071 1633 20105
rect 1583 20047 1633 20071
rect 66187 20105 66237 20129
rect 66187 20071 66195 20105
rect 66229 20071 66237 20105
rect 66187 20047 66237 20071
rect 1583 19769 1633 19793
rect 1583 19735 1591 19769
rect 1625 19735 1633 19769
rect 1583 19711 1633 19735
rect 66187 19769 66237 19793
rect 66187 19735 66195 19769
rect 66229 19735 66237 19769
rect 66187 19711 66237 19735
rect 1583 19433 1633 19457
rect 1583 19399 1591 19433
rect 1625 19399 1633 19433
rect 1583 19375 1633 19399
rect 66187 19433 66237 19457
rect 66187 19399 66195 19433
rect 66229 19399 66237 19433
rect 66187 19375 66237 19399
rect 1583 19097 1633 19121
rect 1583 19063 1591 19097
rect 1625 19063 1633 19097
rect 1583 19039 1633 19063
rect 66187 19097 66237 19121
rect 66187 19063 66195 19097
rect 66229 19063 66237 19097
rect 66187 19039 66237 19063
rect 1583 18761 1633 18785
rect 1583 18727 1591 18761
rect 1625 18727 1633 18761
rect 1583 18703 1633 18727
rect 66187 18761 66237 18785
rect 66187 18727 66195 18761
rect 66229 18727 66237 18761
rect 66187 18703 66237 18727
rect 1583 18425 1633 18449
rect 1583 18391 1591 18425
rect 1625 18391 1633 18425
rect 1583 18367 1633 18391
rect 66187 18425 66237 18449
rect 66187 18391 66195 18425
rect 66229 18391 66237 18425
rect 66187 18367 66237 18391
rect 1583 18089 1633 18113
rect 1583 18055 1591 18089
rect 1625 18055 1633 18089
rect 1583 18031 1633 18055
rect 66187 18089 66237 18113
rect 66187 18055 66195 18089
rect 66229 18055 66237 18089
rect 66187 18031 66237 18055
rect 1583 17753 1633 17777
rect 1583 17719 1591 17753
rect 1625 17719 1633 17753
rect 1583 17695 1633 17719
rect 66187 17753 66237 17777
rect 66187 17719 66195 17753
rect 66229 17719 66237 17753
rect 66187 17695 66237 17719
rect 1583 17417 1633 17441
rect 1583 17383 1591 17417
rect 1625 17383 1633 17417
rect 1583 17359 1633 17383
rect 66187 17417 66237 17441
rect 66187 17383 66195 17417
rect 66229 17383 66237 17417
rect 66187 17359 66237 17383
rect 1583 17081 1633 17105
rect 1583 17047 1591 17081
rect 1625 17047 1633 17081
rect 1583 17023 1633 17047
rect 66187 17081 66237 17105
rect 66187 17047 66195 17081
rect 66229 17047 66237 17081
rect 66187 17023 66237 17047
rect 1583 16745 1633 16769
rect 1583 16711 1591 16745
rect 1625 16711 1633 16745
rect 1583 16687 1633 16711
rect 66187 16745 66237 16769
rect 66187 16711 66195 16745
rect 66229 16711 66237 16745
rect 66187 16687 66237 16711
rect 1583 16409 1633 16433
rect 1583 16375 1591 16409
rect 1625 16375 1633 16409
rect 1583 16351 1633 16375
rect 66187 16409 66237 16433
rect 66187 16375 66195 16409
rect 66229 16375 66237 16409
rect 66187 16351 66237 16375
rect 1583 16073 1633 16097
rect 1583 16039 1591 16073
rect 1625 16039 1633 16073
rect 1583 16015 1633 16039
rect 66187 16073 66237 16097
rect 66187 16039 66195 16073
rect 66229 16039 66237 16073
rect 66187 16015 66237 16039
rect 1583 15737 1633 15761
rect 1583 15703 1591 15737
rect 1625 15703 1633 15737
rect 1583 15679 1633 15703
rect 66187 15737 66237 15761
rect 66187 15703 66195 15737
rect 66229 15703 66237 15737
rect 66187 15679 66237 15703
rect 1583 15401 1633 15425
rect 1583 15367 1591 15401
rect 1625 15367 1633 15401
rect 1583 15343 1633 15367
rect 66187 15401 66237 15425
rect 66187 15367 66195 15401
rect 66229 15367 66237 15401
rect 66187 15343 66237 15367
rect 1583 15065 1633 15089
rect 1583 15031 1591 15065
rect 1625 15031 1633 15065
rect 1583 15007 1633 15031
rect 66187 15065 66237 15089
rect 66187 15031 66195 15065
rect 66229 15031 66237 15065
rect 66187 15007 66237 15031
rect 1583 14729 1633 14753
rect 1583 14695 1591 14729
rect 1625 14695 1633 14729
rect 1583 14671 1633 14695
rect 66187 14729 66237 14753
rect 66187 14695 66195 14729
rect 66229 14695 66237 14729
rect 66187 14671 66237 14695
rect 1583 14393 1633 14417
rect 1583 14359 1591 14393
rect 1625 14359 1633 14393
rect 1583 14335 1633 14359
rect 66187 14393 66237 14417
rect 66187 14359 66195 14393
rect 66229 14359 66237 14393
rect 66187 14335 66237 14359
rect 1583 14057 1633 14081
rect 1583 14023 1591 14057
rect 1625 14023 1633 14057
rect 1583 13999 1633 14023
rect 66187 14057 66237 14081
rect 66187 14023 66195 14057
rect 66229 14023 66237 14057
rect 66187 13999 66237 14023
rect 1583 13721 1633 13745
rect 1583 13687 1591 13721
rect 1625 13687 1633 13721
rect 1583 13663 1633 13687
rect 66187 13721 66237 13745
rect 66187 13687 66195 13721
rect 66229 13687 66237 13721
rect 66187 13663 66237 13687
rect 1583 13385 1633 13409
rect 1583 13351 1591 13385
rect 1625 13351 1633 13385
rect 1583 13327 1633 13351
rect 66187 13385 66237 13409
rect 66187 13351 66195 13385
rect 66229 13351 66237 13385
rect 66187 13327 66237 13351
rect 1583 13049 1633 13073
rect 1583 13015 1591 13049
rect 1625 13015 1633 13049
rect 1583 12991 1633 13015
rect 66187 13049 66237 13073
rect 66187 13015 66195 13049
rect 66229 13015 66237 13049
rect 66187 12991 66237 13015
rect 1583 12713 1633 12737
rect 1583 12679 1591 12713
rect 1625 12679 1633 12713
rect 1583 12655 1633 12679
rect 66187 12713 66237 12737
rect 66187 12679 66195 12713
rect 66229 12679 66237 12713
rect 66187 12655 66237 12679
rect 1583 12377 1633 12401
rect 1583 12343 1591 12377
rect 1625 12343 1633 12377
rect 1583 12319 1633 12343
rect 66187 12377 66237 12401
rect 66187 12343 66195 12377
rect 66229 12343 66237 12377
rect 66187 12319 66237 12343
rect 1583 12041 1633 12065
rect 1583 12007 1591 12041
rect 1625 12007 1633 12041
rect 1583 11983 1633 12007
rect 66187 12041 66237 12065
rect 66187 12007 66195 12041
rect 66229 12007 66237 12041
rect 66187 11983 66237 12007
rect 1583 11705 1633 11729
rect 1583 11671 1591 11705
rect 1625 11671 1633 11705
rect 1583 11647 1633 11671
rect 66187 11705 66237 11729
rect 66187 11671 66195 11705
rect 66229 11671 66237 11705
rect 66187 11647 66237 11671
rect 1583 11369 1633 11393
rect 1583 11335 1591 11369
rect 1625 11335 1633 11369
rect 1583 11311 1633 11335
rect 66187 11369 66237 11393
rect 66187 11335 66195 11369
rect 66229 11335 66237 11369
rect 66187 11311 66237 11335
rect 1583 11033 1633 11057
rect 1583 10999 1591 11033
rect 1625 10999 1633 11033
rect 1583 10975 1633 10999
rect 66187 11033 66237 11057
rect 66187 10999 66195 11033
rect 66229 10999 66237 11033
rect 66187 10975 66237 10999
rect 1583 10697 1633 10721
rect 1583 10663 1591 10697
rect 1625 10663 1633 10697
rect 1583 10639 1633 10663
rect 66187 10697 66237 10721
rect 66187 10663 66195 10697
rect 66229 10663 66237 10697
rect 66187 10639 66237 10663
rect 1583 10361 1633 10385
rect 1583 10327 1591 10361
rect 1625 10327 1633 10361
rect 1583 10303 1633 10327
rect 66187 10361 66237 10385
rect 66187 10327 66195 10361
rect 66229 10327 66237 10361
rect 66187 10303 66237 10327
rect 1583 10025 1633 10049
rect 1583 9991 1591 10025
rect 1625 9991 1633 10025
rect 1583 9967 1633 9991
rect 66187 10025 66237 10049
rect 66187 9991 66195 10025
rect 66229 9991 66237 10025
rect 66187 9967 66237 9991
rect 1583 9689 1633 9713
rect 1583 9655 1591 9689
rect 1625 9655 1633 9689
rect 1583 9631 1633 9655
rect 66187 9689 66237 9713
rect 66187 9655 66195 9689
rect 66229 9655 66237 9689
rect 66187 9631 66237 9655
rect 1583 9353 1633 9377
rect 1583 9319 1591 9353
rect 1625 9319 1633 9353
rect 1583 9295 1633 9319
rect 66187 9353 66237 9377
rect 66187 9319 66195 9353
rect 66229 9319 66237 9353
rect 66187 9295 66237 9319
rect 1583 9017 1633 9041
rect 1583 8983 1591 9017
rect 1625 8983 1633 9017
rect 1583 8959 1633 8983
rect 66187 9017 66237 9041
rect 66187 8983 66195 9017
rect 66229 8983 66237 9017
rect 66187 8959 66237 8983
rect 1583 8681 1633 8705
rect 1583 8647 1591 8681
rect 1625 8647 1633 8681
rect 1583 8623 1633 8647
rect 66187 8681 66237 8705
rect 66187 8647 66195 8681
rect 66229 8647 66237 8681
rect 66187 8623 66237 8647
rect 1583 8345 1633 8369
rect 1583 8311 1591 8345
rect 1625 8311 1633 8345
rect 1583 8287 1633 8311
rect 66187 8345 66237 8369
rect 66187 8311 66195 8345
rect 66229 8311 66237 8345
rect 66187 8287 66237 8311
rect 1583 8009 1633 8033
rect 1583 7975 1591 8009
rect 1625 7975 1633 8009
rect 1583 7951 1633 7975
rect 66187 8009 66237 8033
rect 66187 7975 66195 8009
rect 66229 7975 66237 8009
rect 66187 7951 66237 7975
rect 1583 7673 1633 7697
rect 1583 7639 1591 7673
rect 1625 7639 1633 7673
rect 1583 7615 1633 7639
rect 66187 7673 66237 7697
rect 66187 7639 66195 7673
rect 66229 7639 66237 7673
rect 66187 7615 66237 7639
rect 1583 7337 1633 7361
rect 1583 7303 1591 7337
rect 1625 7303 1633 7337
rect 1583 7279 1633 7303
rect 66187 7337 66237 7361
rect 66187 7303 66195 7337
rect 66229 7303 66237 7337
rect 66187 7279 66237 7303
rect 1583 7001 1633 7025
rect 1583 6967 1591 7001
rect 1625 6967 1633 7001
rect 1583 6943 1633 6967
rect 66187 7001 66237 7025
rect 66187 6967 66195 7001
rect 66229 6967 66237 7001
rect 66187 6943 66237 6967
rect 1583 6665 1633 6689
rect 1583 6631 1591 6665
rect 1625 6631 1633 6665
rect 1583 6607 1633 6631
rect 66187 6665 66237 6689
rect 66187 6631 66195 6665
rect 66229 6631 66237 6665
rect 66187 6607 66237 6631
rect 1583 6329 1633 6353
rect 1583 6295 1591 6329
rect 1625 6295 1633 6329
rect 1583 6271 1633 6295
rect 66187 6329 66237 6353
rect 66187 6295 66195 6329
rect 66229 6295 66237 6329
rect 66187 6271 66237 6295
rect 1583 5993 1633 6017
rect 1583 5959 1591 5993
rect 1625 5959 1633 5993
rect 1583 5935 1633 5959
rect 66187 5993 66237 6017
rect 66187 5959 66195 5993
rect 66229 5959 66237 5993
rect 66187 5935 66237 5959
rect 1583 5657 1633 5681
rect 1583 5623 1591 5657
rect 1625 5623 1633 5657
rect 1583 5599 1633 5623
rect 66187 5657 66237 5681
rect 66187 5623 66195 5657
rect 66229 5623 66237 5657
rect 66187 5599 66237 5623
rect 1583 5321 1633 5345
rect 1583 5287 1591 5321
rect 1625 5287 1633 5321
rect 1583 5263 1633 5287
rect 66187 5321 66237 5345
rect 66187 5287 66195 5321
rect 66229 5287 66237 5321
rect 66187 5263 66237 5287
rect 1583 4985 1633 5009
rect 1583 4951 1591 4985
rect 1625 4951 1633 4985
rect 1583 4927 1633 4951
rect 66187 4985 66237 5009
rect 66187 4951 66195 4985
rect 66229 4951 66237 4985
rect 66187 4927 66237 4951
rect 1583 4649 1633 4673
rect 1583 4615 1591 4649
rect 1625 4615 1633 4649
rect 1583 4591 1633 4615
rect 66187 4649 66237 4673
rect 66187 4615 66195 4649
rect 66229 4615 66237 4649
rect 66187 4591 66237 4615
rect 1583 4313 1633 4337
rect 1583 4279 1591 4313
rect 1625 4279 1633 4313
rect 1583 4255 1633 4279
rect 66187 4313 66237 4337
rect 66187 4279 66195 4313
rect 66229 4279 66237 4313
rect 66187 4255 66237 4279
rect 1583 3977 1633 4001
rect 1583 3943 1591 3977
rect 1625 3943 1633 3977
rect 1583 3919 1633 3943
rect 66187 3977 66237 4001
rect 66187 3943 66195 3977
rect 66229 3943 66237 3977
rect 66187 3919 66237 3943
rect 1583 3641 1633 3665
rect 1583 3607 1591 3641
rect 1625 3607 1633 3641
rect 1583 3583 1633 3607
rect 66187 3641 66237 3665
rect 66187 3607 66195 3641
rect 66229 3607 66237 3641
rect 66187 3583 66237 3607
rect 1583 3305 1633 3329
rect 1583 3271 1591 3305
rect 1625 3271 1633 3305
rect 1583 3247 1633 3271
rect 66187 3305 66237 3329
rect 66187 3271 66195 3305
rect 66229 3271 66237 3305
rect 66187 3247 66237 3271
rect 1583 2969 1633 2993
rect 1583 2935 1591 2969
rect 1625 2935 1633 2969
rect 1583 2911 1633 2935
rect 66187 2969 66237 2993
rect 66187 2935 66195 2969
rect 66229 2935 66237 2969
rect 66187 2911 66237 2935
rect 1583 2633 1633 2657
rect 1583 2599 1591 2633
rect 1625 2599 1633 2633
rect 1583 2575 1633 2599
rect 66187 2633 66237 2657
rect 66187 2599 66195 2633
rect 66229 2599 66237 2633
rect 66187 2575 66237 2599
rect 1583 2297 1633 2321
rect 1583 2263 1591 2297
rect 1625 2263 1633 2297
rect 1583 2239 1633 2263
rect 66187 2297 66237 2321
rect 66187 2263 66195 2297
rect 66229 2263 66237 2297
rect 66187 2239 66237 2263
rect 1583 1961 1633 1985
rect 1583 1927 1591 1961
rect 1625 1927 1633 1961
rect 1583 1903 1633 1927
rect 66187 1961 66237 1985
rect 66187 1927 66195 1961
rect 66229 1927 66237 1961
rect 66187 1903 66237 1927
rect 1919 1625 1969 1649
rect 1919 1591 1927 1625
rect 1961 1591 1969 1625
rect 1919 1567 1969 1591
rect 2255 1625 2305 1649
rect 2255 1591 2263 1625
rect 2297 1591 2305 1625
rect 2255 1567 2305 1591
rect 2591 1625 2641 1649
rect 2591 1591 2599 1625
rect 2633 1591 2641 1625
rect 2591 1567 2641 1591
rect 2927 1625 2977 1649
rect 2927 1591 2935 1625
rect 2969 1591 2977 1625
rect 2927 1567 2977 1591
rect 3263 1625 3313 1649
rect 3263 1591 3271 1625
rect 3305 1591 3313 1625
rect 3263 1567 3313 1591
rect 3599 1625 3649 1649
rect 3599 1591 3607 1625
rect 3641 1591 3649 1625
rect 3599 1567 3649 1591
rect 3935 1625 3985 1649
rect 3935 1591 3943 1625
rect 3977 1591 3985 1625
rect 3935 1567 3985 1591
rect 4271 1625 4321 1649
rect 4271 1591 4279 1625
rect 4313 1591 4321 1625
rect 4271 1567 4321 1591
rect 4607 1625 4657 1649
rect 4607 1591 4615 1625
rect 4649 1591 4657 1625
rect 4607 1567 4657 1591
rect 4943 1625 4993 1649
rect 4943 1591 4951 1625
rect 4985 1591 4993 1625
rect 4943 1567 4993 1591
rect 5279 1625 5329 1649
rect 5279 1591 5287 1625
rect 5321 1591 5329 1625
rect 5279 1567 5329 1591
rect 5615 1625 5665 1649
rect 5615 1591 5623 1625
rect 5657 1591 5665 1625
rect 5615 1567 5665 1591
rect 5951 1625 6001 1649
rect 5951 1591 5959 1625
rect 5993 1591 6001 1625
rect 5951 1567 6001 1591
rect 6287 1625 6337 1649
rect 6287 1591 6295 1625
rect 6329 1591 6337 1625
rect 6287 1567 6337 1591
rect 6623 1625 6673 1649
rect 6623 1591 6631 1625
rect 6665 1591 6673 1625
rect 6623 1567 6673 1591
rect 6959 1625 7009 1649
rect 6959 1591 6967 1625
rect 7001 1591 7009 1625
rect 6959 1567 7009 1591
rect 7295 1625 7345 1649
rect 7295 1591 7303 1625
rect 7337 1591 7345 1625
rect 7295 1567 7345 1591
rect 7631 1625 7681 1649
rect 7631 1591 7639 1625
rect 7673 1591 7681 1625
rect 7631 1567 7681 1591
rect 7967 1625 8017 1649
rect 7967 1591 7975 1625
rect 8009 1591 8017 1625
rect 7967 1567 8017 1591
rect 8303 1625 8353 1649
rect 8303 1591 8311 1625
rect 8345 1591 8353 1625
rect 8303 1567 8353 1591
rect 8639 1625 8689 1649
rect 8639 1591 8647 1625
rect 8681 1591 8689 1625
rect 8639 1567 8689 1591
rect 8975 1625 9025 1649
rect 8975 1591 8983 1625
rect 9017 1591 9025 1625
rect 8975 1567 9025 1591
rect 9311 1625 9361 1649
rect 9311 1591 9319 1625
rect 9353 1591 9361 1625
rect 9311 1567 9361 1591
rect 9647 1625 9697 1649
rect 9647 1591 9655 1625
rect 9689 1591 9697 1625
rect 9647 1567 9697 1591
rect 9983 1625 10033 1649
rect 9983 1591 9991 1625
rect 10025 1591 10033 1625
rect 9983 1567 10033 1591
rect 10319 1625 10369 1649
rect 10319 1591 10327 1625
rect 10361 1591 10369 1625
rect 10319 1567 10369 1591
rect 10655 1625 10705 1649
rect 10655 1591 10663 1625
rect 10697 1591 10705 1625
rect 10655 1567 10705 1591
rect 10991 1625 11041 1649
rect 10991 1591 10999 1625
rect 11033 1591 11041 1625
rect 10991 1567 11041 1591
rect 11327 1625 11377 1649
rect 11327 1591 11335 1625
rect 11369 1591 11377 1625
rect 11327 1567 11377 1591
rect 11663 1625 11713 1649
rect 11663 1591 11671 1625
rect 11705 1591 11713 1625
rect 11663 1567 11713 1591
rect 11999 1625 12049 1649
rect 11999 1591 12007 1625
rect 12041 1591 12049 1625
rect 11999 1567 12049 1591
rect 12335 1625 12385 1649
rect 12335 1591 12343 1625
rect 12377 1591 12385 1625
rect 12335 1567 12385 1591
rect 12671 1625 12721 1649
rect 12671 1591 12679 1625
rect 12713 1591 12721 1625
rect 12671 1567 12721 1591
rect 13007 1625 13057 1649
rect 13007 1591 13015 1625
rect 13049 1591 13057 1625
rect 13007 1567 13057 1591
rect 13343 1625 13393 1649
rect 13343 1591 13351 1625
rect 13385 1591 13393 1625
rect 13343 1567 13393 1591
rect 13679 1625 13729 1649
rect 13679 1591 13687 1625
rect 13721 1591 13729 1625
rect 13679 1567 13729 1591
rect 14015 1625 14065 1649
rect 14015 1591 14023 1625
rect 14057 1591 14065 1625
rect 14015 1567 14065 1591
rect 14351 1625 14401 1649
rect 14351 1591 14359 1625
rect 14393 1591 14401 1625
rect 14351 1567 14401 1591
rect 14687 1625 14737 1649
rect 14687 1591 14695 1625
rect 14729 1591 14737 1625
rect 14687 1567 14737 1591
rect 15023 1625 15073 1649
rect 15023 1591 15031 1625
rect 15065 1591 15073 1625
rect 15023 1567 15073 1591
rect 15359 1625 15409 1649
rect 15359 1591 15367 1625
rect 15401 1591 15409 1625
rect 15359 1567 15409 1591
rect 15695 1625 15745 1649
rect 15695 1591 15703 1625
rect 15737 1591 15745 1625
rect 15695 1567 15745 1591
rect 16031 1625 16081 1649
rect 16031 1591 16039 1625
rect 16073 1591 16081 1625
rect 16031 1567 16081 1591
rect 16367 1625 16417 1649
rect 16367 1591 16375 1625
rect 16409 1591 16417 1625
rect 16367 1567 16417 1591
rect 16703 1625 16753 1649
rect 16703 1591 16711 1625
rect 16745 1591 16753 1625
rect 16703 1567 16753 1591
rect 17039 1625 17089 1649
rect 17039 1591 17047 1625
rect 17081 1591 17089 1625
rect 17039 1567 17089 1591
rect 17375 1625 17425 1649
rect 17375 1591 17383 1625
rect 17417 1591 17425 1625
rect 17375 1567 17425 1591
rect 17711 1625 17761 1649
rect 17711 1591 17719 1625
rect 17753 1591 17761 1625
rect 17711 1567 17761 1591
rect 18047 1625 18097 1649
rect 18047 1591 18055 1625
rect 18089 1591 18097 1625
rect 18047 1567 18097 1591
rect 18383 1625 18433 1649
rect 18383 1591 18391 1625
rect 18425 1591 18433 1625
rect 18383 1567 18433 1591
rect 18719 1625 18769 1649
rect 18719 1591 18727 1625
rect 18761 1591 18769 1625
rect 18719 1567 18769 1591
rect 19055 1625 19105 1649
rect 19055 1591 19063 1625
rect 19097 1591 19105 1625
rect 19055 1567 19105 1591
rect 19391 1625 19441 1649
rect 19391 1591 19399 1625
rect 19433 1591 19441 1625
rect 19391 1567 19441 1591
rect 19727 1625 19777 1649
rect 19727 1591 19735 1625
rect 19769 1591 19777 1625
rect 19727 1567 19777 1591
rect 20063 1625 20113 1649
rect 20063 1591 20071 1625
rect 20105 1591 20113 1625
rect 20063 1567 20113 1591
rect 20399 1625 20449 1649
rect 20399 1591 20407 1625
rect 20441 1591 20449 1625
rect 20399 1567 20449 1591
rect 20735 1625 20785 1649
rect 20735 1591 20743 1625
rect 20777 1591 20785 1625
rect 20735 1567 20785 1591
rect 21071 1625 21121 1649
rect 21071 1591 21079 1625
rect 21113 1591 21121 1625
rect 21071 1567 21121 1591
rect 21407 1625 21457 1649
rect 21407 1591 21415 1625
rect 21449 1591 21457 1625
rect 21407 1567 21457 1591
rect 21743 1625 21793 1649
rect 21743 1591 21751 1625
rect 21785 1591 21793 1625
rect 21743 1567 21793 1591
rect 22079 1625 22129 1649
rect 22079 1591 22087 1625
rect 22121 1591 22129 1625
rect 22079 1567 22129 1591
rect 22415 1625 22465 1649
rect 22415 1591 22423 1625
rect 22457 1591 22465 1625
rect 22415 1567 22465 1591
rect 22751 1625 22801 1649
rect 22751 1591 22759 1625
rect 22793 1591 22801 1625
rect 22751 1567 22801 1591
rect 23087 1625 23137 1649
rect 23087 1591 23095 1625
rect 23129 1591 23137 1625
rect 23087 1567 23137 1591
rect 23423 1625 23473 1649
rect 23423 1591 23431 1625
rect 23465 1591 23473 1625
rect 23423 1567 23473 1591
rect 23759 1625 23809 1649
rect 23759 1591 23767 1625
rect 23801 1591 23809 1625
rect 23759 1567 23809 1591
rect 24095 1625 24145 1649
rect 24095 1591 24103 1625
rect 24137 1591 24145 1625
rect 24095 1567 24145 1591
rect 24431 1625 24481 1649
rect 24431 1591 24439 1625
rect 24473 1591 24481 1625
rect 24431 1567 24481 1591
rect 24767 1625 24817 1649
rect 24767 1591 24775 1625
rect 24809 1591 24817 1625
rect 24767 1567 24817 1591
rect 25103 1625 25153 1649
rect 25103 1591 25111 1625
rect 25145 1591 25153 1625
rect 25103 1567 25153 1591
rect 25439 1625 25489 1649
rect 25439 1591 25447 1625
rect 25481 1591 25489 1625
rect 25439 1567 25489 1591
rect 25775 1625 25825 1649
rect 25775 1591 25783 1625
rect 25817 1591 25825 1625
rect 25775 1567 25825 1591
rect 26111 1625 26161 1649
rect 26111 1591 26119 1625
rect 26153 1591 26161 1625
rect 26111 1567 26161 1591
rect 26447 1625 26497 1649
rect 26447 1591 26455 1625
rect 26489 1591 26497 1625
rect 26447 1567 26497 1591
rect 26783 1625 26833 1649
rect 26783 1591 26791 1625
rect 26825 1591 26833 1625
rect 26783 1567 26833 1591
rect 27119 1625 27169 1649
rect 27119 1591 27127 1625
rect 27161 1591 27169 1625
rect 27119 1567 27169 1591
rect 27455 1625 27505 1649
rect 27455 1591 27463 1625
rect 27497 1591 27505 1625
rect 27455 1567 27505 1591
rect 27791 1625 27841 1649
rect 27791 1591 27799 1625
rect 27833 1591 27841 1625
rect 27791 1567 27841 1591
rect 28127 1625 28177 1649
rect 28127 1591 28135 1625
rect 28169 1591 28177 1625
rect 28127 1567 28177 1591
rect 28463 1625 28513 1649
rect 28463 1591 28471 1625
rect 28505 1591 28513 1625
rect 28463 1567 28513 1591
rect 28799 1625 28849 1649
rect 28799 1591 28807 1625
rect 28841 1591 28849 1625
rect 28799 1567 28849 1591
rect 29135 1625 29185 1649
rect 29135 1591 29143 1625
rect 29177 1591 29185 1625
rect 29135 1567 29185 1591
rect 29471 1625 29521 1649
rect 29471 1591 29479 1625
rect 29513 1591 29521 1625
rect 29471 1567 29521 1591
rect 29807 1625 29857 1649
rect 29807 1591 29815 1625
rect 29849 1591 29857 1625
rect 29807 1567 29857 1591
rect 30143 1625 30193 1649
rect 30143 1591 30151 1625
rect 30185 1591 30193 1625
rect 30143 1567 30193 1591
rect 30479 1625 30529 1649
rect 30479 1591 30487 1625
rect 30521 1591 30529 1625
rect 30479 1567 30529 1591
rect 30815 1625 30865 1649
rect 30815 1591 30823 1625
rect 30857 1591 30865 1625
rect 30815 1567 30865 1591
rect 31151 1625 31201 1649
rect 31151 1591 31159 1625
rect 31193 1591 31201 1625
rect 31151 1567 31201 1591
rect 31487 1625 31537 1649
rect 31487 1591 31495 1625
rect 31529 1591 31537 1625
rect 31487 1567 31537 1591
rect 31823 1625 31873 1649
rect 31823 1591 31831 1625
rect 31865 1591 31873 1625
rect 31823 1567 31873 1591
rect 32159 1625 32209 1649
rect 32159 1591 32167 1625
rect 32201 1591 32209 1625
rect 32159 1567 32209 1591
rect 32495 1625 32545 1649
rect 32495 1591 32503 1625
rect 32537 1591 32545 1625
rect 32495 1567 32545 1591
rect 32831 1625 32881 1649
rect 32831 1591 32839 1625
rect 32873 1591 32881 1625
rect 32831 1567 32881 1591
rect 33167 1625 33217 1649
rect 33167 1591 33175 1625
rect 33209 1591 33217 1625
rect 33167 1567 33217 1591
rect 33503 1625 33553 1649
rect 33503 1591 33511 1625
rect 33545 1591 33553 1625
rect 33503 1567 33553 1591
rect 33839 1625 33889 1649
rect 33839 1591 33847 1625
rect 33881 1591 33889 1625
rect 33839 1567 33889 1591
rect 34175 1625 34225 1649
rect 34175 1591 34183 1625
rect 34217 1591 34225 1625
rect 34175 1567 34225 1591
rect 34511 1625 34561 1649
rect 34511 1591 34519 1625
rect 34553 1591 34561 1625
rect 34511 1567 34561 1591
rect 34847 1625 34897 1649
rect 34847 1591 34855 1625
rect 34889 1591 34897 1625
rect 34847 1567 34897 1591
rect 35183 1625 35233 1649
rect 35183 1591 35191 1625
rect 35225 1591 35233 1625
rect 35183 1567 35233 1591
rect 35519 1625 35569 1649
rect 35519 1591 35527 1625
rect 35561 1591 35569 1625
rect 35519 1567 35569 1591
rect 35855 1625 35905 1649
rect 35855 1591 35863 1625
rect 35897 1591 35905 1625
rect 35855 1567 35905 1591
rect 36191 1625 36241 1649
rect 36191 1591 36199 1625
rect 36233 1591 36241 1625
rect 36191 1567 36241 1591
rect 36527 1625 36577 1649
rect 36527 1591 36535 1625
rect 36569 1591 36577 1625
rect 36527 1567 36577 1591
rect 36863 1625 36913 1649
rect 36863 1591 36871 1625
rect 36905 1591 36913 1625
rect 36863 1567 36913 1591
rect 37199 1625 37249 1649
rect 37199 1591 37207 1625
rect 37241 1591 37249 1625
rect 37199 1567 37249 1591
rect 37535 1625 37585 1649
rect 37535 1591 37543 1625
rect 37577 1591 37585 1625
rect 37535 1567 37585 1591
rect 37871 1625 37921 1649
rect 37871 1591 37879 1625
rect 37913 1591 37921 1625
rect 37871 1567 37921 1591
rect 38207 1625 38257 1649
rect 38207 1591 38215 1625
rect 38249 1591 38257 1625
rect 38207 1567 38257 1591
rect 38543 1625 38593 1649
rect 38543 1591 38551 1625
rect 38585 1591 38593 1625
rect 38543 1567 38593 1591
rect 38879 1625 38929 1649
rect 38879 1591 38887 1625
rect 38921 1591 38929 1625
rect 38879 1567 38929 1591
rect 39215 1625 39265 1649
rect 39215 1591 39223 1625
rect 39257 1591 39265 1625
rect 39215 1567 39265 1591
rect 39551 1625 39601 1649
rect 39551 1591 39559 1625
rect 39593 1591 39601 1625
rect 39551 1567 39601 1591
rect 39887 1625 39937 1649
rect 39887 1591 39895 1625
rect 39929 1591 39937 1625
rect 39887 1567 39937 1591
rect 40223 1625 40273 1649
rect 40223 1591 40231 1625
rect 40265 1591 40273 1625
rect 40223 1567 40273 1591
rect 40559 1625 40609 1649
rect 40559 1591 40567 1625
rect 40601 1591 40609 1625
rect 40559 1567 40609 1591
rect 40895 1625 40945 1649
rect 40895 1591 40903 1625
rect 40937 1591 40945 1625
rect 40895 1567 40945 1591
rect 41231 1625 41281 1649
rect 41231 1591 41239 1625
rect 41273 1591 41281 1625
rect 41231 1567 41281 1591
rect 41567 1625 41617 1649
rect 41567 1591 41575 1625
rect 41609 1591 41617 1625
rect 41567 1567 41617 1591
rect 41903 1625 41953 1649
rect 41903 1591 41911 1625
rect 41945 1591 41953 1625
rect 41903 1567 41953 1591
rect 42239 1625 42289 1649
rect 42239 1591 42247 1625
rect 42281 1591 42289 1625
rect 42239 1567 42289 1591
rect 42575 1625 42625 1649
rect 42575 1591 42583 1625
rect 42617 1591 42625 1625
rect 42575 1567 42625 1591
rect 42911 1625 42961 1649
rect 42911 1591 42919 1625
rect 42953 1591 42961 1625
rect 42911 1567 42961 1591
rect 43247 1625 43297 1649
rect 43247 1591 43255 1625
rect 43289 1591 43297 1625
rect 43247 1567 43297 1591
rect 43583 1625 43633 1649
rect 43583 1591 43591 1625
rect 43625 1591 43633 1625
rect 43583 1567 43633 1591
rect 43919 1625 43969 1649
rect 43919 1591 43927 1625
rect 43961 1591 43969 1625
rect 43919 1567 43969 1591
rect 44255 1625 44305 1649
rect 44255 1591 44263 1625
rect 44297 1591 44305 1625
rect 44255 1567 44305 1591
rect 44591 1625 44641 1649
rect 44591 1591 44599 1625
rect 44633 1591 44641 1625
rect 44591 1567 44641 1591
rect 44927 1625 44977 1649
rect 44927 1591 44935 1625
rect 44969 1591 44977 1625
rect 44927 1567 44977 1591
rect 45263 1625 45313 1649
rect 45263 1591 45271 1625
rect 45305 1591 45313 1625
rect 45263 1567 45313 1591
rect 45599 1625 45649 1649
rect 45599 1591 45607 1625
rect 45641 1591 45649 1625
rect 45599 1567 45649 1591
rect 45935 1625 45985 1649
rect 45935 1591 45943 1625
rect 45977 1591 45985 1625
rect 45935 1567 45985 1591
rect 46271 1625 46321 1649
rect 46271 1591 46279 1625
rect 46313 1591 46321 1625
rect 46271 1567 46321 1591
rect 46607 1625 46657 1649
rect 46607 1591 46615 1625
rect 46649 1591 46657 1625
rect 46607 1567 46657 1591
rect 46943 1625 46993 1649
rect 46943 1591 46951 1625
rect 46985 1591 46993 1625
rect 46943 1567 46993 1591
rect 47279 1625 47329 1649
rect 47279 1591 47287 1625
rect 47321 1591 47329 1625
rect 47279 1567 47329 1591
rect 47615 1625 47665 1649
rect 47615 1591 47623 1625
rect 47657 1591 47665 1625
rect 47615 1567 47665 1591
rect 47951 1625 48001 1649
rect 47951 1591 47959 1625
rect 47993 1591 48001 1625
rect 47951 1567 48001 1591
rect 48287 1625 48337 1649
rect 48287 1591 48295 1625
rect 48329 1591 48337 1625
rect 48287 1567 48337 1591
rect 48623 1625 48673 1649
rect 48623 1591 48631 1625
rect 48665 1591 48673 1625
rect 48623 1567 48673 1591
rect 48959 1625 49009 1649
rect 48959 1591 48967 1625
rect 49001 1591 49009 1625
rect 48959 1567 49009 1591
rect 49295 1625 49345 1649
rect 49295 1591 49303 1625
rect 49337 1591 49345 1625
rect 49295 1567 49345 1591
rect 49631 1625 49681 1649
rect 49631 1591 49639 1625
rect 49673 1591 49681 1625
rect 49631 1567 49681 1591
rect 49967 1625 50017 1649
rect 49967 1591 49975 1625
rect 50009 1591 50017 1625
rect 49967 1567 50017 1591
rect 50303 1625 50353 1649
rect 50303 1591 50311 1625
rect 50345 1591 50353 1625
rect 50303 1567 50353 1591
rect 50639 1625 50689 1649
rect 50639 1591 50647 1625
rect 50681 1591 50689 1625
rect 50639 1567 50689 1591
rect 50975 1625 51025 1649
rect 50975 1591 50983 1625
rect 51017 1591 51025 1625
rect 50975 1567 51025 1591
rect 51311 1625 51361 1649
rect 51311 1591 51319 1625
rect 51353 1591 51361 1625
rect 51311 1567 51361 1591
rect 51647 1625 51697 1649
rect 51647 1591 51655 1625
rect 51689 1591 51697 1625
rect 51647 1567 51697 1591
rect 51983 1625 52033 1649
rect 51983 1591 51991 1625
rect 52025 1591 52033 1625
rect 51983 1567 52033 1591
rect 52319 1625 52369 1649
rect 52319 1591 52327 1625
rect 52361 1591 52369 1625
rect 52319 1567 52369 1591
rect 52655 1625 52705 1649
rect 52655 1591 52663 1625
rect 52697 1591 52705 1625
rect 52655 1567 52705 1591
rect 52991 1625 53041 1649
rect 52991 1591 52999 1625
rect 53033 1591 53041 1625
rect 52991 1567 53041 1591
rect 53327 1625 53377 1649
rect 53327 1591 53335 1625
rect 53369 1591 53377 1625
rect 53327 1567 53377 1591
rect 53663 1625 53713 1649
rect 53663 1591 53671 1625
rect 53705 1591 53713 1625
rect 53663 1567 53713 1591
rect 53999 1625 54049 1649
rect 53999 1591 54007 1625
rect 54041 1591 54049 1625
rect 53999 1567 54049 1591
rect 54335 1625 54385 1649
rect 54335 1591 54343 1625
rect 54377 1591 54385 1625
rect 54335 1567 54385 1591
rect 54671 1625 54721 1649
rect 54671 1591 54679 1625
rect 54713 1591 54721 1625
rect 54671 1567 54721 1591
rect 55007 1625 55057 1649
rect 55007 1591 55015 1625
rect 55049 1591 55057 1625
rect 55007 1567 55057 1591
rect 55343 1625 55393 1649
rect 55343 1591 55351 1625
rect 55385 1591 55393 1625
rect 55343 1567 55393 1591
rect 55679 1625 55729 1649
rect 55679 1591 55687 1625
rect 55721 1591 55729 1625
rect 55679 1567 55729 1591
rect 56015 1625 56065 1649
rect 56015 1591 56023 1625
rect 56057 1591 56065 1625
rect 56015 1567 56065 1591
rect 56351 1625 56401 1649
rect 56351 1591 56359 1625
rect 56393 1591 56401 1625
rect 56351 1567 56401 1591
rect 56687 1625 56737 1649
rect 56687 1591 56695 1625
rect 56729 1591 56737 1625
rect 56687 1567 56737 1591
rect 57023 1625 57073 1649
rect 57023 1591 57031 1625
rect 57065 1591 57073 1625
rect 57023 1567 57073 1591
rect 57359 1625 57409 1649
rect 57359 1591 57367 1625
rect 57401 1591 57409 1625
rect 57359 1567 57409 1591
rect 57695 1625 57745 1649
rect 57695 1591 57703 1625
rect 57737 1591 57745 1625
rect 57695 1567 57745 1591
rect 58031 1625 58081 1649
rect 58031 1591 58039 1625
rect 58073 1591 58081 1625
rect 58031 1567 58081 1591
rect 58367 1625 58417 1649
rect 58367 1591 58375 1625
rect 58409 1591 58417 1625
rect 58367 1567 58417 1591
rect 58703 1625 58753 1649
rect 58703 1591 58711 1625
rect 58745 1591 58753 1625
rect 58703 1567 58753 1591
rect 59039 1625 59089 1649
rect 59039 1591 59047 1625
rect 59081 1591 59089 1625
rect 59039 1567 59089 1591
rect 59375 1625 59425 1649
rect 59375 1591 59383 1625
rect 59417 1591 59425 1625
rect 59375 1567 59425 1591
rect 59711 1625 59761 1649
rect 59711 1591 59719 1625
rect 59753 1591 59761 1625
rect 59711 1567 59761 1591
rect 60047 1625 60097 1649
rect 60047 1591 60055 1625
rect 60089 1591 60097 1625
rect 60047 1567 60097 1591
rect 60383 1625 60433 1649
rect 60383 1591 60391 1625
rect 60425 1591 60433 1625
rect 60383 1567 60433 1591
rect 60719 1625 60769 1649
rect 60719 1591 60727 1625
rect 60761 1591 60769 1625
rect 60719 1567 60769 1591
rect 61055 1625 61105 1649
rect 61055 1591 61063 1625
rect 61097 1591 61105 1625
rect 61055 1567 61105 1591
rect 61391 1625 61441 1649
rect 61391 1591 61399 1625
rect 61433 1591 61441 1625
rect 61391 1567 61441 1591
rect 61727 1625 61777 1649
rect 61727 1591 61735 1625
rect 61769 1591 61777 1625
rect 61727 1567 61777 1591
rect 62063 1625 62113 1649
rect 62063 1591 62071 1625
rect 62105 1591 62113 1625
rect 62063 1567 62113 1591
rect 62399 1625 62449 1649
rect 62399 1591 62407 1625
rect 62441 1591 62449 1625
rect 62399 1567 62449 1591
rect 62735 1625 62785 1649
rect 62735 1591 62743 1625
rect 62777 1591 62785 1625
rect 62735 1567 62785 1591
rect 63071 1625 63121 1649
rect 63071 1591 63079 1625
rect 63113 1591 63121 1625
rect 63071 1567 63121 1591
rect 63407 1625 63457 1649
rect 63407 1591 63415 1625
rect 63449 1591 63457 1625
rect 63407 1567 63457 1591
rect 63743 1625 63793 1649
rect 63743 1591 63751 1625
rect 63785 1591 63793 1625
rect 63743 1567 63793 1591
rect 64079 1625 64129 1649
rect 64079 1591 64087 1625
rect 64121 1591 64129 1625
rect 64079 1567 64129 1591
rect 64415 1625 64465 1649
rect 64415 1591 64423 1625
rect 64457 1591 64465 1625
rect 64415 1567 64465 1591
rect 64751 1625 64801 1649
rect 64751 1591 64759 1625
rect 64793 1591 64801 1625
rect 64751 1567 64801 1591
rect 65087 1625 65137 1649
rect 65087 1591 65095 1625
rect 65129 1591 65137 1625
rect 65087 1567 65137 1591
rect 65423 1625 65473 1649
rect 65423 1591 65431 1625
rect 65465 1591 65473 1625
rect 65423 1567 65473 1591
rect 65759 1625 65809 1649
rect 65759 1591 65767 1625
rect 65801 1591 65809 1625
rect 65759 1567 65809 1591
<< nsubdiffcont >>
rect 1927 51113 1961 51147
rect 2263 51113 2297 51147
rect 2599 51113 2633 51147
rect 2935 51113 2969 51147
rect 3271 51113 3305 51147
rect 3607 51113 3641 51147
rect 3943 51113 3977 51147
rect 4279 51113 4313 51147
rect 4615 51113 4649 51147
rect 4951 51113 4985 51147
rect 5287 51113 5321 51147
rect 5623 51113 5657 51147
rect 5959 51113 5993 51147
rect 6295 51113 6329 51147
rect 6631 51113 6665 51147
rect 6967 51113 7001 51147
rect 7303 51113 7337 51147
rect 7639 51113 7673 51147
rect 7975 51113 8009 51147
rect 8311 51113 8345 51147
rect 8647 51113 8681 51147
rect 8983 51113 9017 51147
rect 9319 51113 9353 51147
rect 9655 51113 9689 51147
rect 9991 51113 10025 51147
rect 10327 51113 10361 51147
rect 10663 51113 10697 51147
rect 10999 51113 11033 51147
rect 11335 51113 11369 51147
rect 11671 51113 11705 51147
rect 12007 51113 12041 51147
rect 12343 51113 12377 51147
rect 12679 51113 12713 51147
rect 13015 51113 13049 51147
rect 13351 51113 13385 51147
rect 13687 51113 13721 51147
rect 14023 51113 14057 51147
rect 14359 51113 14393 51147
rect 14695 51113 14729 51147
rect 15031 51113 15065 51147
rect 15367 51113 15401 51147
rect 15703 51113 15737 51147
rect 16039 51113 16073 51147
rect 16375 51113 16409 51147
rect 16711 51113 16745 51147
rect 17047 51113 17081 51147
rect 17383 51113 17417 51147
rect 17719 51113 17753 51147
rect 18055 51113 18089 51147
rect 18391 51113 18425 51147
rect 18727 51113 18761 51147
rect 19063 51113 19097 51147
rect 19399 51113 19433 51147
rect 19735 51113 19769 51147
rect 20071 51113 20105 51147
rect 20407 51113 20441 51147
rect 20743 51113 20777 51147
rect 21079 51113 21113 51147
rect 21415 51113 21449 51147
rect 21751 51113 21785 51147
rect 22087 51113 22121 51147
rect 22423 51113 22457 51147
rect 22759 51113 22793 51147
rect 23095 51113 23129 51147
rect 23431 51113 23465 51147
rect 23767 51113 23801 51147
rect 24103 51113 24137 51147
rect 24439 51113 24473 51147
rect 24775 51113 24809 51147
rect 25111 51113 25145 51147
rect 25447 51113 25481 51147
rect 25783 51113 25817 51147
rect 26119 51113 26153 51147
rect 26455 51113 26489 51147
rect 26791 51113 26825 51147
rect 27127 51113 27161 51147
rect 27463 51113 27497 51147
rect 27799 51113 27833 51147
rect 28135 51113 28169 51147
rect 28471 51113 28505 51147
rect 28807 51113 28841 51147
rect 29143 51113 29177 51147
rect 29479 51113 29513 51147
rect 29815 51113 29849 51147
rect 30151 51113 30185 51147
rect 30487 51113 30521 51147
rect 30823 51113 30857 51147
rect 31159 51113 31193 51147
rect 31495 51113 31529 51147
rect 31831 51113 31865 51147
rect 32167 51113 32201 51147
rect 32503 51113 32537 51147
rect 32839 51113 32873 51147
rect 33175 51113 33209 51147
rect 33511 51113 33545 51147
rect 33847 51113 33881 51147
rect 34183 51113 34217 51147
rect 34519 51113 34553 51147
rect 34855 51113 34889 51147
rect 35191 51113 35225 51147
rect 35527 51113 35561 51147
rect 35863 51113 35897 51147
rect 36199 51113 36233 51147
rect 36535 51113 36569 51147
rect 36871 51113 36905 51147
rect 37207 51113 37241 51147
rect 37543 51113 37577 51147
rect 37879 51113 37913 51147
rect 38215 51113 38249 51147
rect 38551 51113 38585 51147
rect 38887 51113 38921 51147
rect 39223 51113 39257 51147
rect 39559 51113 39593 51147
rect 39895 51113 39929 51147
rect 40231 51113 40265 51147
rect 40567 51113 40601 51147
rect 40903 51113 40937 51147
rect 41239 51113 41273 51147
rect 41575 51113 41609 51147
rect 41911 51113 41945 51147
rect 42247 51113 42281 51147
rect 42583 51113 42617 51147
rect 42919 51113 42953 51147
rect 43255 51113 43289 51147
rect 43591 51113 43625 51147
rect 43927 51113 43961 51147
rect 44263 51113 44297 51147
rect 44599 51113 44633 51147
rect 44935 51113 44969 51147
rect 45271 51113 45305 51147
rect 45607 51113 45641 51147
rect 45943 51113 45977 51147
rect 46279 51113 46313 51147
rect 46615 51113 46649 51147
rect 46951 51113 46985 51147
rect 47287 51113 47321 51147
rect 47623 51113 47657 51147
rect 47959 51113 47993 51147
rect 48295 51113 48329 51147
rect 48631 51113 48665 51147
rect 48967 51113 49001 51147
rect 49303 51113 49337 51147
rect 49639 51113 49673 51147
rect 49975 51113 50009 51147
rect 50311 51113 50345 51147
rect 50647 51113 50681 51147
rect 50983 51113 51017 51147
rect 51319 51113 51353 51147
rect 51655 51113 51689 51147
rect 51991 51113 52025 51147
rect 52327 51113 52361 51147
rect 52663 51113 52697 51147
rect 52999 51113 53033 51147
rect 53335 51113 53369 51147
rect 53671 51113 53705 51147
rect 54007 51113 54041 51147
rect 54343 51113 54377 51147
rect 54679 51113 54713 51147
rect 55015 51113 55049 51147
rect 55351 51113 55385 51147
rect 55687 51113 55721 51147
rect 56023 51113 56057 51147
rect 56359 51113 56393 51147
rect 56695 51113 56729 51147
rect 57031 51113 57065 51147
rect 57367 51113 57401 51147
rect 57703 51113 57737 51147
rect 58039 51113 58073 51147
rect 58375 51113 58409 51147
rect 58711 51113 58745 51147
rect 59047 51113 59081 51147
rect 59383 51113 59417 51147
rect 59719 51113 59753 51147
rect 60055 51113 60089 51147
rect 60391 51113 60425 51147
rect 60727 51113 60761 51147
rect 61063 51113 61097 51147
rect 61399 51113 61433 51147
rect 61735 51113 61769 51147
rect 62071 51113 62105 51147
rect 62407 51113 62441 51147
rect 62743 51113 62777 51147
rect 63079 51113 63113 51147
rect 63415 51113 63449 51147
rect 63751 51113 63785 51147
rect 64087 51113 64121 51147
rect 64423 51113 64457 51147
rect 64759 51113 64793 51147
rect 65095 51113 65129 51147
rect 65431 51113 65465 51147
rect 65767 51113 65801 51147
rect 1591 50647 1625 50681
rect 66195 50647 66229 50681
rect 1591 50311 1625 50345
rect 66195 50311 66229 50345
rect 1591 49975 1625 50009
rect 66195 49975 66229 50009
rect 1591 49639 1625 49673
rect 66195 49639 66229 49673
rect 1591 49303 1625 49337
rect 66195 49303 66229 49337
rect 1591 48967 1625 49001
rect 66195 48967 66229 49001
rect 1591 48631 1625 48665
rect 66195 48631 66229 48665
rect 1591 48295 1625 48329
rect 66195 48295 66229 48329
rect 1591 47959 1625 47993
rect 66195 47959 66229 47993
rect 1591 47623 1625 47657
rect 66195 47623 66229 47657
rect 1591 47287 1625 47321
rect 66195 47287 66229 47321
rect 1591 46951 1625 46985
rect 66195 46951 66229 46985
rect 1591 46615 1625 46649
rect 66195 46615 66229 46649
rect 1591 46279 1625 46313
rect 66195 46279 66229 46313
rect 1591 45943 1625 45977
rect 66195 45943 66229 45977
rect 1591 45607 1625 45641
rect 66195 45607 66229 45641
rect 1591 45271 1625 45305
rect 66195 45271 66229 45305
rect 1591 44935 1625 44969
rect 66195 44935 66229 44969
rect 1591 44599 1625 44633
rect 66195 44599 66229 44633
rect 1591 44263 1625 44297
rect 66195 44263 66229 44297
rect 1591 43927 1625 43961
rect 66195 43927 66229 43961
rect 1591 43591 1625 43625
rect 66195 43591 66229 43625
rect 1591 43255 1625 43289
rect 66195 43255 66229 43289
rect 1591 42919 1625 42953
rect 66195 42919 66229 42953
rect 1591 42583 1625 42617
rect 66195 42583 66229 42617
rect 1591 42247 1625 42281
rect 66195 42247 66229 42281
rect 1591 41911 1625 41945
rect 66195 41911 66229 41945
rect 1591 41575 1625 41609
rect 66195 41575 66229 41609
rect 1591 41239 1625 41273
rect 66195 41239 66229 41273
rect 1591 40903 1625 40937
rect 66195 40903 66229 40937
rect 1591 40567 1625 40601
rect 66195 40567 66229 40601
rect 1591 40231 1625 40265
rect 66195 40231 66229 40265
rect 1591 39895 1625 39929
rect 66195 39895 66229 39929
rect 1591 39559 1625 39593
rect 66195 39559 66229 39593
rect 1591 39223 1625 39257
rect 66195 39223 66229 39257
rect 1591 38887 1625 38921
rect 66195 38887 66229 38921
rect 1591 38551 1625 38585
rect 66195 38551 66229 38585
rect 1591 38215 1625 38249
rect 66195 38215 66229 38249
rect 1591 37879 1625 37913
rect 66195 37879 66229 37913
rect 1591 37543 1625 37577
rect 66195 37543 66229 37577
rect 1591 37207 1625 37241
rect 66195 37207 66229 37241
rect 1591 36871 1625 36905
rect 66195 36871 66229 36905
rect 1591 36535 1625 36569
rect 66195 36535 66229 36569
rect 1591 36199 1625 36233
rect 66195 36199 66229 36233
rect 1591 35863 1625 35897
rect 66195 35863 66229 35897
rect 1591 35527 1625 35561
rect 66195 35527 66229 35561
rect 1591 35191 1625 35225
rect 66195 35191 66229 35225
rect 1591 34855 1625 34889
rect 66195 34855 66229 34889
rect 1591 34519 1625 34553
rect 66195 34519 66229 34553
rect 1591 34183 1625 34217
rect 66195 34183 66229 34217
rect 1591 33847 1625 33881
rect 66195 33847 66229 33881
rect 1591 33511 1625 33545
rect 66195 33511 66229 33545
rect 1591 33175 1625 33209
rect 66195 33175 66229 33209
rect 1591 32839 1625 32873
rect 66195 32839 66229 32873
rect 1591 32503 1625 32537
rect 66195 32503 66229 32537
rect 1591 32167 1625 32201
rect 66195 32167 66229 32201
rect 1591 31831 1625 31865
rect 66195 31831 66229 31865
rect 1591 31495 1625 31529
rect 66195 31495 66229 31529
rect 1591 31159 1625 31193
rect 66195 31159 66229 31193
rect 1591 30823 1625 30857
rect 66195 30823 66229 30857
rect 1591 30487 1625 30521
rect 66195 30487 66229 30521
rect 1591 30151 1625 30185
rect 66195 30151 66229 30185
rect 1591 29815 1625 29849
rect 66195 29815 66229 29849
rect 1591 29479 1625 29513
rect 66195 29479 66229 29513
rect 1591 29143 1625 29177
rect 66195 29143 66229 29177
rect 1591 28807 1625 28841
rect 66195 28807 66229 28841
rect 1591 28471 1625 28505
rect 66195 28471 66229 28505
rect 1591 28135 1625 28169
rect 66195 28135 66229 28169
rect 1591 27799 1625 27833
rect 66195 27799 66229 27833
rect 1591 27463 1625 27497
rect 66195 27463 66229 27497
rect 1591 27127 1625 27161
rect 66195 27127 66229 27161
rect 1591 26791 1625 26825
rect 66195 26791 66229 26825
rect 1591 26455 1625 26489
rect 66195 26455 66229 26489
rect 1591 26119 1625 26153
rect 66195 26119 66229 26153
rect 1591 25783 1625 25817
rect 66195 25783 66229 25817
rect 1591 25447 1625 25481
rect 66195 25447 66229 25481
rect 1591 25111 1625 25145
rect 66195 25111 66229 25145
rect 1591 24775 1625 24809
rect 66195 24775 66229 24809
rect 1591 24439 1625 24473
rect 66195 24439 66229 24473
rect 1591 24103 1625 24137
rect 66195 24103 66229 24137
rect 1591 23767 1625 23801
rect 66195 23767 66229 23801
rect 1591 23431 1625 23465
rect 66195 23431 66229 23465
rect 1591 23095 1625 23129
rect 66195 23095 66229 23129
rect 1591 22759 1625 22793
rect 66195 22759 66229 22793
rect 1591 22423 1625 22457
rect 66195 22423 66229 22457
rect 1591 22087 1625 22121
rect 66195 22087 66229 22121
rect 1591 21751 1625 21785
rect 66195 21751 66229 21785
rect 1591 21415 1625 21449
rect 66195 21415 66229 21449
rect 1591 21079 1625 21113
rect 66195 21079 66229 21113
rect 1591 20743 1625 20777
rect 66195 20743 66229 20777
rect 1591 20407 1625 20441
rect 66195 20407 66229 20441
rect 1591 20071 1625 20105
rect 66195 20071 66229 20105
rect 1591 19735 1625 19769
rect 66195 19735 66229 19769
rect 1591 19399 1625 19433
rect 66195 19399 66229 19433
rect 1591 19063 1625 19097
rect 66195 19063 66229 19097
rect 1591 18727 1625 18761
rect 66195 18727 66229 18761
rect 1591 18391 1625 18425
rect 66195 18391 66229 18425
rect 1591 18055 1625 18089
rect 66195 18055 66229 18089
rect 1591 17719 1625 17753
rect 66195 17719 66229 17753
rect 1591 17383 1625 17417
rect 66195 17383 66229 17417
rect 1591 17047 1625 17081
rect 66195 17047 66229 17081
rect 1591 16711 1625 16745
rect 66195 16711 66229 16745
rect 1591 16375 1625 16409
rect 66195 16375 66229 16409
rect 1591 16039 1625 16073
rect 66195 16039 66229 16073
rect 1591 15703 1625 15737
rect 66195 15703 66229 15737
rect 1591 15367 1625 15401
rect 66195 15367 66229 15401
rect 1591 15031 1625 15065
rect 66195 15031 66229 15065
rect 1591 14695 1625 14729
rect 66195 14695 66229 14729
rect 1591 14359 1625 14393
rect 66195 14359 66229 14393
rect 1591 14023 1625 14057
rect 66195 14023 66229 14057
rect 1591 13687 1625 13721
rect 66195 13687 66229 13721
rect 1591 13351 1625 13385
rect 66195 13351 66229 13385
rect 1591 13015 1625 13049
rect 66195 13015 66229 13049
rect 1591 12679 1625 12713
rect 66195 12679 66229 12713
rect 1591 12343 1625 12377
rect 66195 12343 66229 12377
rect 1591 12007 1625 12041
rect 66195 12007 66229 12041
rect 1591 11671 1625 11705
rect 66195 11671 66229 11705
rect 1591 11335 1625 11369
rect 66195 11335 66229 11369
rect 1591 10999 1625 11033
rect 66195 10999 66229 11033
rect 1591 10663 1625 10697
rect 66195 10663 66229 10697
rect 1591 10327 1625 10361
rect 66195 10327 66229 10361
rect 1591 9991 1625 10025
rect 66195 9991 66229 10025
rect 1591 9655 1625 9689
rect 66195 9655 66229 9689
rect 1591 9319 1625 9353
rect 66195 9319 66229 9353
rect 1591 8983 1625 9017
rect 66195 8983 66229 9017
rect 1591 8647 1625 8681
rect 66195 8647 66229 8681
rect 1591 8311 1625 8345
rect 66195 8311 66229 8345
rect 1591 7975 1625 8009
rect 66195 7975 66229 8009
rect 1591 7639 1625 7673
rect 66195 7639 66229 7673
rect 1591 7303 1625 7337
rect 66195 7303 66229 7337
rect 1591 6967 1625 7001
rect 66195 6967 66229 7001
rect 1591 6631 1625 6665
rect 66195 6631 66229 6665
rect 1591 6295 1625 6329
rect 66195 6295 66229 6329
rect 1591 5959 1625 5993
rect 66195 5959 66229 5993
rect 1591 5623 1625 5657
rect 66195 5623 66229 5657
rect 1591 5287 1625 5321
rect 66195 5287 66229 5321
rect 1591 4951 1625 4985
rect 66195 4951 66229 4985
rect 1591 4615 1625 4649
rect 66195 4615 66229 4649
rect 1591 4279 1625 4313
rect 66195 4279 66229 4313
rect 1591 3943 1625 3977
rect 66195 3943 66229 3977
rect 1591 3607 1625 3641
rect 66195 3607 66229 3641
rect 1591 3271 1625 3305
rect 66195 3271 66229 3305
rect 1591 2935 1625 2969
rect 66195 2935 66229 2969
rect 1591 2599 1625 2633
rect 66195 2599 66229 2633
rect 1591 2263 1625 2297
rect 66195 2263 66229 2297
rect 1591 1927 1625 1961
rect 66195 1927 66229 1961
rect 1927 1591 1961 1625
rect 2263 1591 2297 1625
rect 2599 1591 2633 1625
rect 2935 1591 2969 1625
rect 3271 1591 3305 1625
rect 3607 1591 3641 1625
rect 3943 1591 3977 1625
rect 4279 1591 4313 1625
rect 4615 1591 4649 1625
rect 4951 1591 4985 1625
rect 5287 1591 5321 1625
rect 5623 1591 5657 1625
rect 5959 1591 5993 1625
rect 6295 1591 6329 1625
rect 6631 1591 6665 1625
rect 6967 1591 7001 1625
rect 7303 1591 7337 1625
rect 7639 1591 7673 1625
rect 7975 1591 8009 1625
rect 8311 1591 8345 1625
rect 8647 1591 8681 1625
rect 8983 1591 9017 1625
rect 9319 1591 9353 1625
rect 9655 1591 9689 1625
rect 9991 1591 10025 1625
rect 10327 1591 10361 1625
rect 10663 1591 10697 1625
rect 10999 1591 11033 1625
rect 11335 1591 11369 1625
rect 11671 1591 11705 1625
rect 12007 1591 12041 1625
rect 12343 1591 12377 1625
rect 12679 1591 12713 1625
rect 13015 1591 13049 1625
rect 13351 1591 13385 1625
rect 13687 1591 13721 1625
rect 14023 1591 14057 1625
rect 14359 1591 14393 1625
rect 14695 1591 14729 1625
rect 15031 1591 15065 1625
rect 15367 1591 15401 1625
rect 15703 1591 15737 1625
rect 16039 1591 16073 1625
rect 16375 1591 16409 1625
rect 16711 1591 16745 1625
rect 17047 1591 17081 1625
rect 17383 1591 17417 1625
rect 17719 1591 17753 1625
rect 18055 1591 18089 1625
rect 18391 1591 18425 1625
rect 18727 1591 18761 1625
rect 19063 1591 19097 1625
rect 19399 1591 19433 1625
rect 19735 1591 19769 1625
rect 20071 1591 20105 1625
rect 20407 1591 20441 1625
rect 20743 1591 20777 1625
rect 21079 1591 21113 1625
rect 21415 1591 21449 1625
rect 21751 1591 21785 1625
rect 22087 1591 22121 1625
rect 22423 1591 22457 1625
rect 22759 1591 22793 1625
rect 23095 1591 23129 1625
rect 23431 1591 23465 1625
rect 23767 1591 23801 1625
rect 24103 1591 24137 1625
rect 24439 1591 24473 1625
rect 24775 1591 24809 1625
rect 25111 1591 25145 1625
rect 25447 1591 25481 1625
rect 25783 1591 25817 1625
rect 26119 1591 26153 1625
rect 26455 1591 26489 1625
rect 26791 1591 26825 1625
rect 27127 1591 27161 1625
rect 27463 1591 27497 1625
rect 27799 1591 27833 1625
rect 28135 1591 28169 1625
rect 28471 1591 28505 1625
rect 28807 1591 28841 1625
rect 29143 1591 29177 1625
rect 29479 1591 29513 1625
rect 29815 1591 29849 1625
rect 30151 1591 30185 1625
rect 30487 1591 30521 1625
rect 30823 1591 30857 1625
rect 31159 1591 31193 1625
rect 31495 1591 31529 1625
rect 31831 1591 31865 1625
rect 32167 1591 32201 1625
rect 32503 1591 32537 1625
rect 32839 1591 32873 1625
rect 33175 1591 33209 1625
rect 33511 1591 33545 1625
rect 33847 1591 33881 1625
rect 34183 1591 34217 1625
rect 34519 1591 34553 1625
rect 34855 1591 34889 1625
rect 35191 1591 35225 1625
rect 35527 1591 35561 1625
rect 35863 1591 35897 1625
rect 36199 1591 36233 1625
rect 36535 1591 36569 1625
rect 36871 1591 36905 1625
rect 37207 1591 37241 1625
rect 37543 1591 37577 1625
rect 37879 1591 37913 1625
rect 38215 1591 38249 1625
rect 38551 1591 38585 1625
rect 38887 1591 38921 1625
rect 39223 1591 39257 1625
rect 39559 1591 39593 1625
rect 39895 1591 39929 1625
rect 40231 1591 40265 1625
rect 40567 1591 40601 1625
rect 40903 1591 40937 1625
rect 41239 1591 41273 1625
rect 41575 1591 41609 1625
rect 41911 1591 41945 1625
rect 42247 1591 42281 1625
rect 42583 1591 42617 1625
rect 42919 1591 42953 1625
rect 43255 1591 43289 1625
rect 43591 1591 43625 1625
rect 43927 1591 43961 1625
rect 44263 1591 44297 1625
rect 44599 1591 44633 1625
rect 44935 1591 44969 1625
rect 45271 1591 45305 1625
rect 45607 1591 45641 1625
rect 45943 1591 45977 1625
rect 46279 1591 46313 1625
rect 46615 1591 46649 1625
rect 46951 1591 46985 1625
rect 47287 1591 47321 1625
rect 47623 1591 47657 1625
rect 47959 1591 47993 1625
rect 48295 1591 48329 1625
rect 48631 1591 48665 1625
rect 48967 1591 49001 1625
rect 49303 1591 49337 1625
rect 49639 1591 49673 1625
rect 49975 1591 50009 1625
rect 50311 1591 50345 1625
rect 50647 1591 50681 1625
rect 50983 1591 51017 1625
rect 51319 1591 51353 1625
rect 51655 1591 51689 1625
rect 51991 1591 52025 1625
rect 52327 1591 52361 1625
rect 52663 1591 52697 1625
rect 52999 1591 53033 1625
rect 53335 1591 53369 1625
rect 53671 1591 53705 1625
rect 54007 1591 54041 1625
rect 54343 1591 54377 1625
rect 54679 1591 54713 1625
rect 55015 1591 55049 1625
rect 55351 1591 55385 1625
rect 55687 1591 55721 1625
rect 56023 1591 56057 1625
rect 56359 1591 56393 1625
rect 56695 1591 56729 1625
rect 57031 1591 57065 1625
rect 57367 1591 57401 1625
rect 57703 1591 57737 1625
rect 58039 1591 58073 1625
rect 58375 1591 58409 1625
rect 58711 1591 58745 1625
rect 59047 1591 59081 1625
rect 59383 1591 59417 1625
rect 59719 1591 59753 1625
rect 60055 1591 60089 1625
rect 60391 1591 60425 1625
rect 60727 1591 60761 1625
rect 61063 1591 61097 1625
rect 61399 1591 61433 1625
rect 61735 1591 61769 1625
rect 62071 1591 62105 1625
rect 62407 1591 62441 1625
rect 62743 1591 62777 1625
rect 63079 1591 63113 1625
rect 63415 1591 63449 1625
rect 63751 1591 63785 1625
rect 64087 1591 64121 1625
rect 64423 1591 64457 1625
rect 64759 1591 64793 1625
rect 65095 1591 65129 1625
rect 65431 1591 65465 1625
rect 65767 1591 65801 1625
<< locali >>
rect 1927 51147 1961 51163
rect 1927 51097 1961 51113
rect 2263 51147 2297 51163
rect 2263 51097 2297 51113
rect 2599 51147 2633 51163
rect 2599 51097 2633 51113
rect 2935 51147 2969 51163
rect 2935 51097 2969 51113
rect 3271 51147 3305 51163
rect 3271 51097 3305 51113
rect 3607 51147 3641 51163
rect 3607 51097 3641 51113
rect 3943 51147 3977 51163
rect 3943 51097 3977 51113
rect 4279 51147 4313 51163
rect 4279 51097 4313 51113
rect 4615 51147 4649 51163
rect 4615 51097 4649 51113
rect 4951 51147 4985 51163
rect 4951 51097 4985 51113
rect 5287 51147 5321 51163
rect 5287 51097 5321 51113
rect 5623 51147 5657 51163
rect 5623 51097 5657 51113
rect 5959 51147 5993 51163
rect 5959 51097 5993 51113
rect 6295 51147 6329 51163
rect 6295 51097 6329 51113
rect 6631 51147 6665 51163
rect 6631 51097 6665 51113
rect 6967 51147 7001 51163
rect 6967 51097 7001 51113
rect 7303 51147 7337 51163
rect 7303 51097 7337 51113
rect 7639 51147 7673 51163
rect 7639 51097 7673 51113
rect 7975 51147 8009 51163
rect 7975 51097 8009 51113
rect 8311 51147 8345 51163
rect 8311 51097 8345 51113
rect 8647 51147 8681 51163
rect 8647 51097 8681 51113
rect 8983 51147 9017 51163
rect 8983 51097 9017 51113
rect 9319 51147 9353 51163
rect 9319 51097 9353 51113
rect 9655 51147 9689 51163
rect 9655 51097 9689 51113
rect 9991 51147 10025 51163
rect 9991 51097 10025 51113
rect 10327 51147 10361 51163
rect 10327 51097 10361 51113
rect 10663 51147 10697 51163
rect 10663 51097 10697 51113
rect 10999 51147 11033 51163
rect 10999 51097 11033 51113
rect 11335 51147 11369 51163
rect 11335 51097 11369 51113
rect 11671 51147 11705 51163
rect 11671 51097 11705 51113
rect 12007 51147 12041 51163
rect 12007 51097 12041 51113
rect 12343 51147 12377 51163
rect 12343 51097 12377 51113
rect 12679 51147 12713 51163
rect 12679 51097 12713 51113
rect 13015 51147 13049 51163
rect 13015 51097 13049 51113
rect 13351 51147 13385 51163
rect 13351 51097 13385 51113
rect 13687 51147 13721 51163
rect 13687 51097 13721 51113
rect 14023 51147 14057 51163
rect 14023 51097 14057 51113
rect 14359 51147 14393 51163
rect 14359 51097 14393 51113
rect 14695 51147 14729 51163
rect 14695 51097 14729 51113
rect 15031 51147 15065 51163
rect 15031 51097 15065 51113
rect 15367 51147 15401 51163
rect 15367 51097 15401 51113
rect 15703 51147 15737 51163
rect 15703 51097 15737 51113
rect 16039 51147 16073 51163
rect 16039 51097 16073 51113
rect 16375 51147 16409 51163
rect 16375 51097 16409 51113
rect 16711 51147 16745 51163
rect 16711 51097 16745 51113
rect 17047 51147 17081 51163
rect 17047 51097 17081 51113
rect 17383 51147 17417 51163
rect 17383 51097 17417 51113
rect 17719 51147 17753 51163
rect 17719 51097 17753 51113
rect 18055 51147 18089 51163
rect 18055 51097 18089 51113
rect 18391 51147 18425 51163
rect 18391 51097 18425 51113
rect 18727 51147 18761 51163
rect 18727 51097 18761 51113
rect 19063 51147 19097 51163
rect 19063 51097 19097 51113
rect 19399 51147 19433 51163
rect 19399 51097 19433 51113
rect 19735 51147 19769 51163
rect 19735 51097 19769 51113
rect 20071 51147 20105 51163
rect 20071 51097 20105 51113
rect 20407 51147 20441 51163
rect 20407 51097 20441 51113
rect 20743 51147 20777 51163
rect 20743 51097 20777 51113
rect 21079 51147 21113 51163
rect 21079 51097 21113 51113
rect 21415 51147 21449 51163
rect 21415 51097 21449 51113
rect 21751 51147 21785 51163
rect 21751 51097 21785 51113
rect 22087 51147 22121 51163
rect 22087 51097 22121 51113
rect 22423 51147 22457 51163
rect 22423 51097 22457 51113
rect 22759 51147 22793 51163
rect 22759 51097 22793 51113
rect 23095 51147 23129 51163
rect 23095 51097 23129 51113
rect 23431 51147 23465 51163
rect 23431 51097 23465 51113
rect 23767 51147 23801 51163
rect 23767 51097 23801 51113
rect 24103 51147 24137 51163
rect 24103 51097 24137 51113
rect 24439 51147 24473 51163
rect 24439 51097 24473 51113
rect 24775 51147 24809 51163
rect 24775 51097 24809 51113
rect 25111 51147 25145 51163
rect 25111 51097 25145 51113
rect 25447 51147 25481 51163
rect 25447 51097 25481 51113
rect 25783 51147 25817 51163
rect 25783 51097 25817 51113
rect 26119 51147 26153 51163
rect 26119 51097 26153 51113
rect 26455 51147 26489 51163
rect 26455 51097 26489 51113
rect 26791 51147 26825 51163
rect 26791 51097 26825 51113
rect 27127 51147 27161 51163
rect 27127 51097 27161 51113
rect 27463 51147 27497 51163
rect 27463 51097 27497 51113
rect 27799 51147 27833 51163
rect 27799 51097 27833 51113
rect 28135 51147 28169 51163
rect 28135 51097 28169 51113
rect 28471 51147 28505 51163
rect 28471 51097 28505 51113
rect 28807 51147 28841 51163
rect 28807 51097 28841 51113
rect 29143 51147 29177 51163
rect 29143 51097 29177 51113
rect 29479 51147 29513 51163
rect 29479 51097 29513 51113
rect 29815 51147 29849 51163
rect 29815 51097 29849 51113
rect 30151 51147 30185 51163
rect 30151 51097 30185 51113
rect 30487 51147 30521 51163
rect 30487 51097 30521 51113
rect 30823 51147 30857 51163
rect 30823 51097 30857 51113
rect 31159 51147 31193 51163
rect 31159 51097 31193 51113
rect 31495 51147 31529 51163
rect 31495 51097 31529 51113
rect 31831 51147 31865 51163
rect 31831 51097 31865 51113
rect 32167 51147 32201 51163
rect 32167 51097 32201 51113
rect 32503 51147 32537 51163
rect 32503 51097 32537 51113
rect 32839 51147 32873 51163
rect 32839 51097 32873 51113
rect 33175 51147 33209 51163
rect 33175 51097 33209 51113
rect 33511 51147 33545 51163
rect 33511 51097 33545 51113
rect 33847 51147 33881 51163
rect 33847 51097 33881 51113
rect 34183 51147 34217 51163
rect 34183 51097 34217 51113
rect 34519 51147 34553 51163
rect 34519 51097 34553 51113
rect 34855 51147 34889 51163
rect 34855 51097 34889 51113
rect 35191 51147 35225 51163
rect 35191 51097 35225 51113
rect 35527 51147 35561 51163
rect 35527 51097 35561 51113
rect 35863 51147 35897 51163
rect 35863 51097 35897 51113
rect 36199 51147 36233 51163
rect 36199 51097 36233 51113
rect 36535 51147 36569 51163
rect 36535 51097 36569 51113
rect 36871 51147 36905 51163
rect 36871 51097 36905 51113
rect 37207 51147 37241 51163
rect 37207 51097 37241 51113
rect 37543 51147 37577 51163
rect 37543 51097 37577 51113
rect 37879 51147 37913 51163
rect 37879 51097 37913 51113
rect 38215 51147 38249 51163
rect 38215 51097 38249 51113
rect 38551 51147 38585 51163
rect 38551 51097 38585 51113
rect 38887 51147 38921 51163
rect 38887 51097 38921 51113
rect 39223 51147 39257 51163
rect 39223 51097 39257 51113
rect 39559 51147 39593 51163
rect 39559 51097 39593 51113
rect 39895 51147 39929 51163
rect 39895 51097 39929 51113
rect 40231 51147 40265 51163
rect 40231 51097 40265 51113
rect 40567 51147 40601 51163
rect 40567 51097 40601 51113
rect 40903 51147 40937 51163
rect 40903 51097 40937 51113
rect 41239 51147 41273 51163
rect 41239 51097 41273 51113
rect 41575 51147 41609 51163
rect 41575 51097 41609 51113
rect 41911 51147 41945 51163
rect 41911 51097 41945 51113
rect 42247 51147 42281 51163
rect 42247 51097 42281 51113
rect 42583 51147 42617 51163
rect 42583 51097 42617 51113
rect 42919 51147 42953 51163
rect 42919 51097 42953 51113
rect 43255 51147 43289 51163
rect 43255 51097 43289 51113
rect 43591 51147 43625 51163
rect 43591 51097 43625 51113
rect 43927 51147 43961 51163
rect 43927 51097 43961 51113
rect 44263 51147 44297 51163
rect 44263 51097 44297 51113
rect 44599 51147 44633 51163
rect 44599 51097 44633 51113
rect 44935 51147 44969 51163
rect 44935 51097 44969 51113
rect 45271 51147 45305 51163
rect 45271 51097 45305 51113
rect 45607 51147 45641 51163
rect 45607 51097 45641 51113
rect 45943 51147 45977 51163
rect 45943 51097 45977 51113
rect 46279 51147 46313 51163
rect 46279 51097 46313 51113
rect 46615 51147 46649 51163
rect 46615 51097 46649 51113
rect 46951 51147 46985 51163
rect 46951 51097 46985 51113
rect 47287 51147 47321 51163
rect 47287 51097 47321 51113
rect 47623 51147 47657 51163
rect 47623 51097 47657 51113
rect 47959 51147 47993 51163
rect 47959 51097 47993 51113
rect 48295 51147 48329 51163
rect 48295 51097 48329 51113
rect 48631 51147 48665 51163
rect 48631 51097 48665 51113
rect 48967 51147 49001 51163
rect 48967 51097 49001 51113
rect 49303 51147 49337 51163
rect 49303 51097 49337 51113
rect 49639 51147 49673 51163
rect 49639 51097 49673 51113
rect 49975 51147 50009 51163
rect 49975 51097 50009 51113
rect 50311 51147 50345 51163
rect 50311 51097 50345 51113
rect 50647 51147 50681 51163
rect 50647 51097 50681 51113
rect 50983 51147 51017 51163
rect 50983 51097 51017 51113
rect 51319 51147 51353 51163
rect 51319 51097 51353 51113
rect 51655 51147 51689 51163
rect 51655 51097 51689 51113
rect 51991 51147 52025 51163
rect 51991 51097 52025 51113
rect 52327 51147 52361 51163
rect 52327 51097 52361 51113
rect 52663 51147 52697 51163
rect 52663 51097 52697 51113
rect 52999 51147 53033 51163
rect 52999 51097 53033 51113
rect 53335 51147 53369 51163
rect 53335 51097 53369 51113
rect 53671 51147 53705 51163
rect 53671 51097 53705 51113
rect 54007 51147 54041 51163
rect 54007 51097 54041 51113
rect 54343 51147 54377 51163
rect 54343 51097 54377 51113
rect 54679 51147 54713 51163
rect 54679 51097 54713 51113
rect 55015 51147 55049 51163
rect 55015 51097 55049 51113
rect 55351 51147 55385 51163
rect 55351 51097 55385 51113
rect 55687 51147 55721 51163
rect 55687 51097 55721 51113
rect 56023 51147 56057 51163
rect 56023 51097 56057 51113
rect 56359 51147 56393 51163
rect 56359 51097 56393 51113
rect 56695 51147 56729 51163
rect 56695 51097 56729 51113
rect 57031 51147 57065 51163
rect 57031 51097 57065 51113
rect 57367 51147 57401 51163
rect 57367 51097 57401 51113
rect 57703 51147 57737 51163
rect 57703 51097 57737 51113
rect 58039 51147 58073 51163
rect 58039 51097 58073 51113
rect 58375 51147 58409 51163
rect 58375 51097 58409 51113
rect 58711 51147 58745 51163
rect 58711 51097 58745 51113
rect 59047 51147 59081 51163
rect 59047 51097 59081 51113
rect 59383 51147 59417 51163
rect 59383 51097 59417 51113
rect 59719 51147 59753 51163
rect 59719 51097 59753 51113
rect 60055 51147 60089 51163
rect 60055 51097 60089 51113
rect 60391 51147 60425 51163
rect 60391 51097 60425 51113
rect 60727 51147 60761 51163
rect 60727 51097 60761 51113
rect 61063 51147 61097 51163
rect 61063 51097 61097 51113
rect 61399 51147 61433 51163
rect 61399 51097 61433 51113
rect 61735 51147 61769 51163
rect 61735 51097 61769 51113
rect 62071 51147 62105 51163
rect 62071 51097 62105 51113
rect 62407 51147 62441 51163
rect 62407 51097 62441 51113
rect 62743 51147 62777 51163
rect 62743 51097 62777 51113
rect 63079 51147 63113 51163
rect 63079 51097 63113 51113
rect 63415 51147 63449 51163
rect 63415 51097 63449 51113
rect 63751 51147 63785 51163
rect 63751 51097 63785 51113
rect 64087 51147 64121 51163
rect 64087 51097 64121 51113
rect 64423 51147 64457 51163
rect 64423 51097 64457 51113
rect 64759 51147 64793 51163
rect 64759 51097 64793 51113
rect 65095 51147 65129 51163
rect 65095 51097 65129 51113
rect 65431 51147 65465 51163
rect 65431 51097 65465 51113
rect 65767 51147 65801 51163
rect 65767 51097 65801 51113
rect 1591 50681 1625 50697
rect 1591 50631 1625 50647
rect 66195 50681 66229 50697
rect 66195 50631 66229 50647
rect 1591 50345 1625 50361
rect 1591 50295 1625 50311
rect 66195 50345 66229 50361
rect 66195 50295 66229 50311
rect 1591 50009 1625 50025
rect 1591 49959 1625 49975
rect 66195 50009 66229 50025
rect 66195 49959 66229 49975
rect 1591 49673 1625 49689
rect 1591 49623 1625 49639
rect 66195 49673 66229 49689
rect 66195 49623 66229 49639
rect 1591 49337 1625 49353
rect 1591 49287 1625 49303
rect 66195 49337 66229 49353
rect 66195 49287 66229 49303
rect 1591 49001 1625 49017
rect 1591 48951 1625 48967
rect 66195 49001 66229 49017
rect 66195 48951 66229 48967
rect 1591 48665 1625 48681
rect 1591 48615 1625 48631
rect 66195 48665 66229 48681
rect 66195 48615 66229 48631
rect 1591 48329 1625 48345
rect 1591 48279 1625 48295
rect 66195 48329 66229 48345
rect 66195 48279 66229 48295
rect 1591 47993 1625 48009
rect 1591 47943 1625 47959
rect 66195 47993 66229 48009
rect 66195 47943 66229 47959
rect 1591 47657 1625 47673
rect 1591 47607 1625 47623
rect 66195 47657 66229 47673
rect 66195 47607 66229 47623
rect 1591 47321 1625 47337
rect 1591 47271 1625 47287
rect 66195 47321 66229 47337
rect 66195 47271 66229 47287
rect 1591 46985 1625 47001
rect 1591 46935 1625 46951
rect 66195 46985 66229 47001
rect 66195 46935 66229 46951
rect 1591 46649 1625 46665
rect 1591 46599 1625 46615
rect 66195 46649 66229 46665
rect 66195 46599 66229 46615
rect 1591 46313 1625 46329
rect 1591 46263 1625 46279
rect 66195 46313 66229 46329
rect 66195 46263 66229 46279
rect 1591 45977 1625 45993
rect 1591 45927 1625 45943
rect 66195 45977 66229 45993
rect 66195 45927 66229 45943
rect 1591 45641 1625 45657
rect 1591 45591 1625 45607
rect 66195 45641 66229 45657
rect 66195 45591 66229 45607
rect 1591 45305 1625 45321
rect 1591 45255 1625 45271
rect 66195 45305 66229 45321
rect 66195 45255 66229 45271
rect 1591 44969 1625 44985
rect 1591 44919 1625 44935
rect 66195 44969 66229 44985
rect 66195 44919 66229 44935
rect 1591 44633 1625 44649
rect 1591 44583 1625 44599
rect 66195 44633 66229 44649
rect 66195 44583 66229 44599
rect 1591 44297 1625 44313
rect 1591 44247 1625 44263
rect 66195 44297 66229 44313
rect 66195 44247 66229 44263
rect 1591 43961 1625 43977
rect 1591 43911 1625 43927
rect 66195 43961 66229 43977
rect 66195 43911 66229 43927
rect 1591 43625 1625 43641
rect 1591 43575 1625 43591
rect 66195 43625 66229 43641
rect 66195 43575 66229 43591
rect 1591 43289 1625 43305
rect 1591 43239 1625 43255
rect 66195 43289 66229 43305
rect 66195 43239 66229 43255
rect 1591 42953 1625 42969
rect 1591 42903 1625 42919
rect 66195 42953 66229 42969
rect 66195 42903 66229 42919
rect 1591 42617 1625 42633
rect 1591 42567 1625 42583
rect 66195 42617 66229 42633
rect 66195 42567 66229 42583
rect 1591 42281 1625 42297
rect 1591 42231 1625 42247
rect 66195 42281 66229 42297
rect 66195 42231 66229 42247
rect 1591 41945 1625 41961
rect 1591 41895 1625 41911
rect 66195 41945 66229 41961
rect 66195 41895 66229 41911
rect 1591 41609 1625 41625
rect 1591 41559 1625 41575
rect 66195 41609 66229 41625
rect 66195 41559 66229 41575
rect 1591 41273 1625 41289
rect 1591 41223 1625 41239
rect 66195 41273 66229 41289
rect 66195 41223 66229 41239
rect 1591 40937 1625 40953
rect 1591 40887 1625 40903
rect 66195 40937 66229 40953
rect 66195 40887 66229 40903
rect 1591 40601 1625 40617
rect 1591 40551 1625 40567
rect 66195 40601 66229 40617
rect 66195 40551 66229 40567
rect 1591 40265 1625 40281
rect 1591 40215 1625 40231
rect 66195 40265 66229 40281
rect 66195 40215 66229 40231
rect 1591 39929 1625 39945
rect 1591 39879 1625 39895
rect 66195 39929 66229 39945
rect 66195 39879 66229 39895
rect 1591 39593 1625 39609
rect 1591 39543 1625 39559
rect 66195 39593 66229 39609
rect 66195 39543 66229 39559
rect 1591 39257 1625 39273
rect 1591 39207 1625 39223
rect 66195 39257 66229 39273
rect 66195 39207 66229 39223
rect 1591 38921 1625 38937
rect 1591 38871 1625 38887
rect 66195 38921 66229 38937
rect 66195 38871 66229 38887
rect 1591 38585 1625 38601
rect 1591 38535 1625 38551
rect 66195 38585 66229 38601
rect 66195 38535 66229 38551
rect 1591 38249 1625 38265
rect 1591 38199 1625 38215
rect 66195 38249 66229 38265
rect 66195 38199 66229 38215
rect 1591 37913 1625 37929
rect 1591 37863 1625 37879
rect 66195 37913 66229 37929
rect 66195 37863 66229 37879
rect 1591 37577 1625 37593
rect 1591 37527 1625 37543
rect 66195 37577 66229 37593
rect 66195 37527 66229 37543
rect 1591 37241 1625 37257
rect 1591 37191 1625 37207
rect 66195 37241 66229 37257
rect 66195 37191 66229 37207
rect 1591 36905 1625 36921
rect 1591 36855 1625 36871
rect 66195 36905 66229 36921
rect 66195 36855 66229 36871
rect 1591 36569 1625 36585
rect 1591 36519 1625 36535
rect 66195 36569 66229 36585
rect 66195 36519 66229 36535
rect 1591 36233 1625 36249
rect 1591 36183 1625 36199
rect 66195 36233 66229 36249
rect 66195 36183 66229 36199
rect 1591 35897 1625 35913
rect 1591 35847 1625 35863
rect 66195 35897 66229 35913
rect 66195 35847 66229 35863
rect 1591 35561 1625 35577
rect 1591 35511 1625 35527
rect 66195 35561 66229 35577
rect 66195 35511 66229 35527
rect 1591 35225 1625 35241
rect 1591 35175 1625 35191
rect 66195 35225 66229 35241
rect 66195 35175 66229 35191
rect 1591 34889 1625 34905
rect 1591 34839 1625 34855
rect 66195 34889 66229 34905
rect 66195 34839 66229 34855
rect 1591 34553 1625 34569
rect 1591 34503 1625 34519
rect 66195 34553 66229 34569
rect 66195 34503 66229 34519
rect 1591 34217 1625 34233
rect 1591 34167 1625 34183
rect 66195 34217 66229 34233
rect 66195 34167 66229 34183
rect 1591 33881 1625 33897
rect 1591 33831 1625 33847
rect 66195 33881 66229 33897
rect 66195 33831 66229 33847
rect 1591 33545 1625 33561
rect 1591 33495 1625 33511
rect 66195 33545 66229 33561
rect 66195 33495 66229 33511
rect 1591 33209 1625 33225
rect 1591 33159 1625 33175
rect 66195 33209 66229 33225
rect 66195 33159 66229 33175
rect 1591 32873 1625 32889
rect 1591 32823 1625 32839
rect 66195 32873 66229 32889
rect 66195 32823 66229 32839
rect 1591 32537 1625 32553
rect 1591 32487 1625 32503
rect 66195 32537 66229 32553
rect 66195 32487 66229 32503
rect 1591 32201 1625 32217
rect 1591 32151 1625 32167
rect 66195 32201 66229 32217
rect 66195 32151 66229 32167
rect 1591 31865 1625 31881
rect 1591 31815 1625 31831
rect 66195 31865 66229 31881
rect 66195 31815 66229 31831
rect 1591 31529 1625 31545
rect 1591 31479 1625 31495
rect 66195 31529 66229 31545
rect 66195 31479 66229 31495
rect 1591 31193 1625 31209
rect 1591 31143 1625 31159
rect 66195 31193 66229 31209
rect 66195 31143 66229 31159
rect 1591 30857 1625 30873
rect 1591 30807 1625 30823
rect 66195 30857 66229 30873
rect 66195 30807 66229 30823
rect 1591 30521 1625 30537
rect 1591 30471 1625 30487
rect 66195 30521 66229 30537
rect 66195 30471 66229 30487
rect 1591 30185 1625 30201
rect 1591 30135 1625 30151
rect 66195 30185 66229 30201
rect 66195 30135 66229 30151
rect 1591 29849 1625 29865
rect 1591 29799 1625 29815
rect 66195 29849 66229 29865
rect 66195 29799 66229 29815
rect 1591 29513 1625 29529
rect 1591 29463 1625 29479
rect 66195 29513 66229 29529
rect 66195 29463 66229 29479
rect 1591 29177 1625 29193
rect 1591 29127 1625 29143
rect 66195 29177 66229 29193
rect 66195 29127 66229 29143
rect 1591 28841 1625 28857
rect 1591 28791 1625 28807
rect 66195 28841 66229 28857
rect 66195 28791 66229 28807
rect 1591 28505 1625 28521
rect 1591 28455 1625 28471
rect 66195 28505 66229 28521
rect 66195 28455 66229 28471
rect 1591 28169 1625 28185
rect 1591 28119 1625 28135
rect 66195 28169 66229 28185
rect 66195 28119 66229 28135
rect 1591 27833 1625 27849
rect 1591 27783 1625 27799
rect 66195 27833 66229 27849
rect 66195 27783 66229 27799
rect 1591 27497 1625 27513
rect 1591 27447 1625 27463
rect 66195 27497 66229 27513
rect 66195 27447 66229 27463
rect 1591 27161 1625 27177
rect 1591 27111 1625 27127
rect 66195 27161 66229 27177
rect 66195 27111 66229 27127
rect 1591 26825 1625 26841
rect 1591 26775 1625 26791
rect 66195 26825 66229 26841
rect 66195 26775 66229 26791
rect 1591 26489 1625 26505
rect 1591 26439 1625 26455
rect 66195 26489 66229 26505
rect 66195 26439 66229 26455
rect 1591 26153 1625 26169
rect 1591 26103 1625 26119
rect 66195 26153 66229 26169
rect 66195 26103 66229 26119
rect 1591 25817 1625 25833
rect 1591 25767 1625 25783
rect 66195 25817 66229 25833
rect 66195 25767 66229 25783
rect 1591 25481 1625 25497
rect 1591 25431 1625 25447
rect 66195 25481 66229 25497
rect 66195 25431 66229 25447
rect 1591 25145 1625 25161
rect 1591 25095 1625 25111
rect 66195 25145 66229 25161
rect 66195 25095 66229 25111
rect 1591 24809 1625 24825
rect 1591 24759 1625 24775
rect 66195 24809 66229 24825
rect 66195 24759 66229 24775
rect 1591 24473 1625 24489
rect 1591 24423 1625 24439
rect 66195 24473 66229 24489
rect 66195 24423 66229 24439
rect 1591 24137 1625 24153
rect 1591 24087 1625 24103
rect 66195 24137 66229 24153
rect 66195 24087 66229 24103
rect 1591 23801 1625 23817
rect 1591 23751 1625 23767
rect 66195 23801 66229 23817
rect 66195 23751 66229 23767
rect 1591 23465 1625 23481
rect 1591 23415 1625 23431
rect 66195 23465 66229 23481
rect 66195 23415 66229 23431
rect 1591 23129 1625 23145
rect 1591 23079 1625 23095
rect 66195 23129 66229 23145
rect 66195 23079 66229 23095
rect 1591 22793 1625 22809
rect 1591 22743 1625 22759
rect 66195 22793 66229 22809
rect 66195 22743 66229 22759
rect 1591 22457 1625 22473
rect 1591 22407 1625 22423
rect 66195 22457 66229 22473
rect 66195 22407 66229 22423
rect 1591 22121 1625 22137
rect 1591 22071 1625 22087
rect 66195 22121 66229 22137
rect 66195 22071 66229 22087
rect 1591 21785 1625 21801
rect 1591 21735 1625 21751
rect 66195 21785 66229 21801
rect 66195 21735 66229 21751
rect 1591 21449 1625 21465
rect 1591 21399 1625 21415
rect 66195 21449 66229 21465
rect 66195 21399 66229 21415
rect 1591 21113 1625 21129
rect 1591 21063 1625 21079
rect 66195 21113 66229 21129
rect 66195 21063 66229 21079
rect 1591 20777 1625 20793
rect 1591 20727 1625 20743
rect 66195 20777 66229 20793
rect 66195 20727 66229 20743
rect 1591 20441 1625 20457
rect 1591 20391 1625 20407
rect 66195 20441 66229 20457
rect 66195 20391 66229 20407
rect 1591 20105 1625 20121
rect 1591 20055 1625 20071
rect 66195 20105 66229 20121
rect 66195 20055 66229 20071
rect 1591 19769 1625 19785
rect 1591 19719 1625 19735
rect 66195 19769 66229 19785
rect 66195 19719 66229 19735
rect 1591 19433 1625 19449
rect 1591 19383 1625 19399
rect 66195 19433 66229 19449
rect 66195 19383 66229 19399
rect 1591 19097 1625 19113
rect 1591 19047 1625 19063
rect 66195 19097 66229 19113
rect 66195 19047 66229 19063
rect 1591 18761 1625 18777
rect 1591 18711 1625 18727
rect 66195 18761 66229 18777
rect 66195 18711 66229 18727
rect 1591 18425 1625 18441
rect 1591 18375 1625 18391
rect 66195 18425 66229 18441
rect 66195 18375 66229 18391
rect 1591 18089 1625 18105
rect 1591 18039 1625 18055
rect 66195 18089 66229 18105
rect 66195 18039 66229 18055
rect 1591 17753 1625 17769
rect 1591 17703 1625 17719
rect 66195 17753 66229 17769
rect 66195 17703 66229 17719
rect 1591 17417 1625 17433
rect 1591 17367 1625 17383
rect 66195 17417 66229 17433
rect 66195 17367 66229 17383
rect 1591 17081 1625 17097
rect 1591 17031 1625 17047
rect 66195 17081 66229 17097
rect 66195 17031 66229 17047
rect 1591 16745 1625 16761
rect 1591 16695 1625 16711
rect 66195 16745 66229 16761
rect 66195 16695 66229 16711
rect 1591 16409 1625 16425
rect 1591 16359 1625 16375
rect 66195 16409 66229 16425
rect 66195 16359 66229 16375
rect 1591 16073 1625 16089
rect 1591 16023 1625 16039
rect 66195 16073 66229 16089
rect 66195 16023 66229 16039
rect 1591 15737 1625 15753
rect 1591 15687 1625 15703
rect 66195 15737 66229 15753
rect 66195 15687 66229 15703
rect 1591 15401 1625 15417
rect 1591 15351 1625 15367
rect 66195 15401 66229 15417
rect 66195 15351 66229 15367
rect 1591 15065 1625 15081
rect 1591 15015 1625 15031
rect 66195 15065 66229 15081
rect 66195 15015 66229 15031
rect 1591 14729 1625 14745
rect 1591 14679 1625 14695
rect 66195 14729 66229 14745
rect 66195 14679 66229 14695
rect 1591 14393 1625 14409
rect 1591 14343 1625 14359
rect 66195 14393 66229 14409
rect 66195 14343 66229 14359
rect 1591 14057 1625 14073
rect 1591 14007 1625 14023
rect 66195 14057 66229 14073
rect 66195 14007 66229 14023
rect 1591 13721 1625 13737
rect 1591 13671 1625 13687
rect 66195 13721 66229 13737
rect 66195 13671 66229 13687
rect 1591 13385 1625 13401
rect 1591 13335 1625 13351
rect 66195 13385 66229 13401
rect 66195 13335 66229 13351
rect 1591 13049 1625 13065
rect 1591 12999 1625 13015
rect 66195 13049 66229 13065
rect 66195 12999 66229 13015
rect 1591 12713 1625 12729
rect 1591 12663 1625 12679
rect 66195 12713 66229 12729
rect 66195 12663 66229 12679
rect 1591 12377 1625 12393
rect 1591 12327 1625 12343
rect 66195 12377 66229 12393
rect 66195 12327 66229 12343
rect 1591 12041 1625 12057
rect 1591 11991 1625 12007
rect 66195 12041 66229 12057
rect 66195 11991 66229 12007
rect 1591 11705 1625 11721
rect 1591 11655 1625 11671
rect 66195 11705 66229 11721
rect 66195 11655 66229 11671
rect 1591 11369 1625 11385
rect 1591 11319 1625 11335
rect 66195 11369 66229 11385
rect 66195 11319 66229 11335
rect 1591 11033 1625 11049
rect 1591 10983 1625 10999
rect 66195 11033 66229 11049
rect 66195 10983 66229 10999
rect 1591 10697 1625 10713
rect 1591 10647 1625 10663
rect 66195 10697 66229 10713
rect 66195 10647 66229 10663
rect 1591 10361 1625 10377
rect 1591 10311 1625 10327
rect 66195 10361 66229 10377
rect 66195 10311 66229 10327
rect 1591 10025 1625 10041
rect 1591 9975 1625 9991
rect 66195 10025 66229 10041
rect 66195 9975 66229 9991
rect 1591 9689 1625 9705
rect 1591 9639 1625 9655
rect 66195 9689 66229 9705
rect 66195 9639 66229 9655
rect 1591 9353 1625 9369
rect 1591 9303 1625 9319
rect 66195 9353 66229 9369
rect 66195 9303 66229 9319
rect 1591 9017 1625 9033
rect 1591 8967 1625 8983
rect 66195 9017 66229 9033
rect 66195 8967 66229 8983
rect 1591 8681 1625 8697
rect 1591 8631 1625 8647
rect 66195 8681 66229 8697
rect 66195 8631 66229 8647
rect 1591 8345 1625 8361
rect 1591 8295 1625 8311
rect 66195 8345 66229 8361
rect 66195 8295 66229 8311
rect 1591 8009 1625 8025
rect 1591 7959 1625 7975
rect 66195 8009 66229 8025
rect 66195 7959 66229 7975
rect 1591 7673 1625 7689
rect 1591 7623 1625 7639
rect 66195 7673 66229 7689
rect 66195 7623 66229 7639
rect 1591 7337 1625 7353
rect 1591 7287 1625 7303
rect 66195 7337 66229 7353
rect 66195 7287 66229 7303
rect 1591 7001 1625 7017
rect 1591 6951 1625 6967
rect 66195 7001 66229 7017
rect 66195 6951 66229 6967
rect 1591 6665 1625 6681
rect 1591 6615 1625 6631
rect 66195 6665 66229 6681
rect 66195 6615 66229 6631
rect 1591 6329 1625 6345
rect 1591 6279 1625 6295
rect 66195 6329 66229 6345
rect 66195 6279 66229 6295
rect 1591 5993 1625 6009
rect 1591 5943 1625 5959
rect 66195 5993 66229 6009
rect 66195 5943 66229 5959
rect 1591 5657 1625 5673
rect 1591 5607 1625 5623
rect 66195 5657 66229 5673
rect 66195 5607 66229 5623
rect 1591 5321 1625 5337
rect 1591 5271 1625 5287
rect 66195 5321 66229 5337
rect 66195 5271 66229 5287
rect 1591 4985 1625 5001
rect 1591 4935 1625 4951
rect 66195 4985 66229 5001
rect 66195 4935 66229 4951
rect 1591 4649 1625 4665
rect 1591 4599 1625 4615
rect 66195 4649 66229 4665
rect 66195 4599 66229 4615
rect 1591 4313 1625 4329
rect 1591 4263 1625 4279
rect 66195 4313 66229 4329
rect 66195 4263 66229 4279
rect 1591 3977 1625 3993
rect 1591 3927 1625 3943
rect 66195 3977 66229 3993
rect 66195 3927 66229 3943
rect 1591 3641 1625 3657
rect 1591 3591 1625 3607
rect 66195 3641 66229 3657
rect 66195 3591 66229 3607
rect 1591 3305 1625 3321
rect 1591 3255 1625 3271
rect 66195 3305 66229 3321
rect 66195 3255 66229 3271
rect 1591 2969 1625 2985
rect 1591 2919 1625 2935
rect 66195 2969 66229 2985
rect 66195 2919 66229 2935
rect 1591 2633 1625 2649
rect 1591 2583 1625 2599
rect 66195 2633 66229 2649
rect 66195 2583 66229 2599
rect 1591 2297 1625 2313
rect 1591 2247 1625 2263
rect 66195 2297 66229 2313
rect 66195 2247 66229 2263
rect 1591 1961 1625 1977
rect 1591 1911 1625 1927
rect 66195 1961 66229 1977
rect 66195 1911 66229 1927
rect 1927 1625 1961 1641
rect 1927 1575 1961 1591
rect 2263 1625 2297 1641
rect 2263 1575 2297 1591
rect 2599 1625 2633 1641
rect 2599 1575 2633 1591
rect 2935 1625 2969 1641
rect 2935 1575 2969 1591
rect 3271 1625 3305 1641
rect 3271 1575 3305 1591
rect 3607 1625 3641 1641
rect 3607 1575 3641 1591
rect 3943 1625 3977 1641
rect 3943 1575 3977 1591
rect 4279 1625 4313 1641
rect 4279 1575 4313 1591
rect 4615 1625 4649 1641
rect 4615 1575 4649 1591
rect 4951 1625 4985 1641
rect 4951 1575 4985 1591
rect 5287 1625 5321 1641
rect 5287 1575 5321 1591
rect 5623 1625 5657 1641
rect 5623 1575 5657 1591
rect 5959 1625 5993 1641
rect 5959 1575 5993 1591
rect 6295 1625 6329 1641
rect 6295 1575 6329 1591
rect 6631 1625 6665 1641
rect 6631 1575 6665 1591
rect 6967 1625 7001 1641
rect 6967 1575 7001 1591
rect 7303 1625 7337 1641
rect 7303 1575 7337 1591
rect 7639 1625 7673 1641
rect 7639 1575 7673 1591
rect 7975 1625 8009 1641
rect 7975 1575 8009 1591
rect 8311 1625 8345 1641
rect 8311 1575 8345 1591
rect 8647 1625 8681 1641
rect 8647 1575 8681 1591
rect 8983 1625 9017 1641
rect 8983 1575 9017 1591
rect 9319 1625 9353 1641
rect 9319 1575 9353 1591
rect 9655 1625 9689 1641
rect 9655 1575 9689 1591
rect 9991 1625 10025 1641
rect 9991 1575 10025 1591
rect 10327 1625 10361 1641
rect 10327 1575 10361 1591
rect 10663 1625 10697 1641
rect 10663 1575 10697 1591
rect 10999 1625 11033 1641
rect 10999 1575 11033 1591
rect 11335 1625 11369 1641
rect 11335 1575 11369 1591
rect 11671 1625 11705 1641
rect 11671 1575 11705 1591
rect 12007 1625 12041 1641
rect 12007 1575 12041 1591
rect 12343 1625 12377 1641
rect 12343 1575 12377 1591
rect 12679 1625 12713 1641
rect 12679 1575 12713 1591
rect 13015 1625 13049 1641
rect 13015 1575 13049 1591
rect 13351 1625 13385 1641
rect 13351 1575 13385 1591
rect 13687 1625 13721 1641
rect 13687 1575 13721 1591
rect 14023 1625 14057 1641
rect 14023 1575 14057 1591
rect 14359 1625 14393 1641
rect 14359 1575 14393 1591
rect 14695 1625 14729 1641
rect 14695 1575 14729 1591
rect 15031 1625 15065 1641
rect 15031 1575 15065 1591
rect 15367 1625 15401 1641
rect 15367 1575 15401 1591
rect 15703 1625 15737 1641
rect 15703 1575 15737 1591
rect 16039 1625 16073 1641
rect 16039 1575 16073 1591
rect 16375 1625 16409 1641
rect 16375 1575 16409 1591
rect 16711 1625 16745 1641
rect 16711 1575 16745 1591
rect 17047 1625 17081 1641
rect 17047 1575 17081 1591
rect 17383 1625 17417 1641
rect 17383 1575 17417 1591
rect 17719 1625 17753 1641
rect 17719 1575 17753 1591
rect 18055 1625 18089 1641
rect 18055 1575 18089 1591
rect 18391 1625 18425 1641
rect 18391 1575 18425 1591
rect 18727 1625 18761 1641
rect 18727 1575 18761 1591
rect 19063 1625 19097 1641
rect 19063 1575 19097 1591
rect 19399 1625 19433 1641
rect 19399 1575 19433 1591
rect 19735 1625 19769 1641
rect 19735 1575 19769 1591
rect 20071 1625 20105 1641
rect 20071 1575 20105 1591
rect 20407 1625 20441 1641
rect 20407 1575 20441 1591
rect 20743 1625 20777 1641
rect 20743 1575 20777 1591
rect 21079 1625 21113 1641
rect 21079 1575 21113 1591
rect 21415 1625 21449 1641
rect 21415 1575 21449 1591
rect 21751 1625 21785 1641
rect 21751 1575 21785 1591
rect 22087 1625 22121 1641
rect 22087 1575 22121 1591
rect 22423 1625 22457 1641
rect 22423 1575 22457 1591
rect 22759 1625 22793 1641
rect 22759 1575 22793 1591
rect 23095 1625 23129 1641
rect 23095 1575 23129 1591
rect 23431 1625 23465 1641
rect 23431 1575 23465 1591
rect 23767 1625 23801 1641
rect 23767 1575 23801 1591
rect 24103 1625 24137 1641
rect 24103 1575 24137 1591
rect 24439 1625 24473 1641
rect 24439 1575 24473 1591
rect 24775 1625 24809 1641
rect 24775 1575 24809 1591
rect 25111 1625 25145 1641
rect 25111 1575 25145 1591
rect 25447 1625 25481 1641
rect 25447 1575 25481 1591
rect 25783 1625 25817 1641
rect 25783 1575 25817 1591
rect 26119 1625 26153 1641
rect 26119 1575 26153 1591
rect 26455 1625 26489 1641
rect 26455 1575 26489 1591
rect 26791 1625 26825 1641
rect 26791 1575 26825 1591
rect 27127 1625 27161 1641
rect 27127 1575 27161 1591
rect 27463 1625 27497 1641
rect 27463 1575 27497 1591
rect 27799 1625 27833 1641
rect 27799 1575 27833 1591
rect 28135 1625 28169 1641
rect 28135 1575 28169 1591
rect 28471 1625 28505 1641
rect 28471 1575 28505 1591
rect 28807 1625 28841 1641
rect 28807 1575 28841 1591
rect 29143 1625 29177 1641
rect 29143 1575 29177 1591
rect 29479 1625 29513 1641
rect 29479 1575 29513 1591
rect 29815 1625 29849 1641
rect 29815 1575 29849 1591
rect 30151 1625 30185 1641
rect 30151 1575 30185 1591
rect 30487 1625 30521 1641
rect 30487 1575 30521 1591
rect 30823 1625 30857 1641
rect 30823 1575 30857 1591
rect 31159 1625 31193 1641
rect 31159 1575 31193 1591
rect 31495 1625 31529 1641
rect 31495 1575 31529 1591
rect 31831 1625 31865 1641
rect 31831 1575 31865 1591
rect 32167 1625 32201 1641
rect 32167 1575 32201 1591
rect 32503 1625 32537 1641
rect 32503 1575 32537 1591
rect 32839 1625 32873 1641
rect 32839 1575 32873 1591
rect 33175 1625 33209 1641
rect 33175 1575 33209 1591
rect 33511 1625 33545 1641
rect 33511 1575 33545 1591
rect 33847 1625 33881 1641
rect 33847 1575 33881 1591
rect 34183 1625 34217 1641
rect 34183 1575 34217 1591
rect 34519 1625 34553 1641
rect 34519 1575 34553 1591
rect 34855 1625 34889 1641
rect 34855 1575 34889 1591
rect 35191 1625 35225 1641
rect 35191 1575 35225 1591
rect 35527 1625 35561 1641
rect 35527 1575 35561 1591
rect 35863 1625 35897 1641
rect 35863 1575 35897 1591
rect 36199 1625 36233 1641
rect 36199 1575 36233 1591
rect 36535 1625 36569 1641
rect 36535 1575 36569 1591
rect 36871 1625 36905 1641
rect 36871 1575 36905 1591
rect 37207 1625 37241 1641
rect 37207 1575 37241 1591
rect 37543 1625 37577 1641
rect 37543 1575 37577 1591
rect 37879 1625 37913 1641
rect 37879 1575 37913 1591
rect 38215 1625 38249 1641
rect 38215 1575 38249 1591
rect 38551 1625 38585 1641
rect 38551 1575 38585 1591
rect 38887 1625 38921 1641
rect 38887 1575 38921 1591
rect 39223 1625 39257 1641
rect 39223 1575 39257 1591
rect 39559 1625 39593 1641
rect 39559 1575 39593 1591
rect 39895 1625 39929 1641
rect 39895 1575 39929 1591
rect 40231 1625 40265 1641
rect 40231 1575 40265 1591
rect 40567 1625 40601 1641
rect 40567 1575 40601 1591
rect 40903 1625 40937 1641
rect 40903 1575 40937 1591
rect 41239 1625 41273 1641
rect 41239 1575 41273 1591
rect 41575 1625 41609 1641
rect 41575 1575 41609 1591
rect 41911 1625 41945 1641
rect 41911 1575 41945 1591
rect 42247 1625 42281 1641
rect 42247 1575 42281 1591
rect 42583 1625 42617 1641
rect 42583 1575 42617 1591
rect 42919 1625 42953 1641
rect 42919 1575 42953 1591
rect 43255 1625 43289 1641
rect 43255 1575 43289 1591
rect 43591 1625 43625 1641
rect 43591 1575 43625 1591
rect 43927 1625 43961 1641
rect 43927 1575 43961 1591
rect 44263 1625 44297 1641
rect 44263 1575 44297 1591
rect 44599 1625 44633 1641
rect 44599 1575 44633 1591
rect 44935 1625 44969 1641
rect 44935 1575 44969 1591
rect 45271 1625 45305 1641
rect 45271 1575 45305 1591
rect 45607 1625 45641 1641
rect 45607 1575 45641 1591
rect 45943 1625 45977 1641
rect 45943 1575 45977 1591
rect 46279 1625 46313 1641
rect 46279 1575 46313 1591
rect 46615 1625 46649 1641
rect 46615 1575 46649 1591
rect 46951 1625 46985 1641
rect 46951 1575 46985 1591
rect 47287 1625 47321 1641
rect 47287 1575 47321 1591
rect 47623 1625 47657 1641
rect 47623 1575 47657 1591
rect 47959 1625 47993 1641
rect 47959 1575 47993 1591
rect 48295 1625 48329 1641
rect 48295 1575 48329 1591
rect 48631 1625 48665 1641
rect 48631 1575 48665 1591
rect 48967 1625 49001 1641
rect 48967 1575 49001 1591
rect 49303 1625 49337 1641
rect 49303 1575 49337 1591
rect 49639 1625 49673 1641
rect 49639 1575 49673 1591
rect 49975 1625 50009 1641
rect 49975 1575 50009 1591
rect 50311 1625 50345 1641
rect 50311 1575 50345 1591
rect 50647 1625 50681 1641
rect 50647 1575 50681 1591
rect 50983 1625 51017 1641
rect 50983 1575 51017 1591
rect 51319 1625 51353 1641
rect 51319 1575 51353 1591
rect 51655 1625 51689 1641
rect 51655 1575 51689 1591
rect 51991 1625 52025 1641
rect 51991 1575 52025 1591
rect 52327 1625 52361 1641
rect 52327 1575 52361 1591
rect 52663 1625 52697 1641
rect 52663 1575 52697 1591
rect 52999 1625 53033 1641
rect 52999 1575 53033 1591
rect 53335 1625 53369 1641
rect 53335 1575 53369 1591
rect 53671 1625 53705 1641
rect 53671 1575 53705 1591
rect 54007 1625 54041 1641
rect 54007 1575 54041 1591
rect 54343 1625 54377 1641
rect 54343 1575 54377 1591
rect 54679 1625 54713 1641
rect 54679 1575 54713 1591
rect 55015 1625 55049 1641
rect 55015 1575 55049 1591
rect 55351 1625 55385 1641
rect 55351 1575 55385 1591
rect 55687 1625 55721 1641
rect 55687 1575 55721 1591
rect 56023 1625 56057 1641
rect 56023 1575 56057 1591
rect 56359 1625 56393 1641
rect 56359 1575 56393 1591
rect 56695 1625 56729 1641
rect 56695 1575 56729 1591
rect 57031 1625 57065 1641
rect 57031 1575 57065 1591
rect 57367 1625 57401 1641
rect 57367 1575 57401 1591
rect 57703 1625 57737 1641
rect 57703 1575 57737 1591
rect 58039 1625 58073 1641
rect 58039 1575 58073 1591
rect 58375 1625 58409 1641
rect 58375 1575 58409 1591
rect 58711 1625 58745 1641
rect 58711 1575 58745 1591
rect 59047 1625 59081 1641
rect 59047 1575 59081 1591
rect 59383 1625 59417 1641
rect 59383 1575 59417 1591
rect 59719 1625 59753 1641
rect 59719 1575 59753 1591
rect 60055 1625 60089 1641
rect 60055 1575 60089 1591
rect 60391 1625 60425 1641
rect 60391 1575 60425 1591
rect 60727 1625 60761 1641
rect 60727 1575 60761 1591
rect 61063 1625 61097 1641
rect 61063 1575 61097 1591
rect 61399 1625 61433 1641
rect 61399 1575 61433 1591
rect 61735 1625 61769 1641
rect 61735 1575 61769 1591
rect 62071 1625 62105 1641
rect 62071 1575 62105 1591
rect 62407 1625 62441 1641
rect 62407 1575 62441 1591
rect 62743 1625 62777 1641
rect 62743 1575 62777 1591
rect 63079 1625 63113 1641
rect 63079 1575 63113 1591
rect 63415 1625 63449 1641
rect 63415 1575 63449 1591
rect 63751 1625 63785 1641
rect 63751 1575 63785 1591
rect 64087 1625 64121 1641
rect 64087 1575 64121 1591
rect 64423 1625 64457 1641
rect 64423 1575 64457 1591
rect 64759 1625 64793 1641
rect 64759 1575 64793 1591
rect 65095 1625 65129 1641
rect 65095 1575 65129 1591
rect 65431 1625 65465 1641
rect 65431 1575 65465 1591
rect 65767 1625 65801 1641
rect 65767 1575 65801 1591
<< viali >>
rect 1927 51113 1961 51147
rect 2263 51113 2297 51147
rect 2599 51113 2633 51147
rect 2935 51113 2969 51147
rect 3271 51113 3305 51147
rect 3607 51113 3641 51147
rect 3943 51113 3977 51147
rect 4279 51113 4313 51147
rect 4615 51113 4649 51147
rect 4951 51113 4985 51147
rect 5287 51113 5321 51147
rect 5623 51113 5657 51147
rect 5959 51113 5993 51147
rect 6295 51113 6329 51147
rect 6631 51113 6665 51147
rect 6967 51113 7001 51147
rect 7303 51113 7337 51147
rect 7639 51113 7673 51147
rect 7975 51113 8009 51147
rect 8311 51113 8345 51147
rect 8647 51113 8681 51147
rect 8983 51113 9017 51147
rect 9319 51113 9353 51147
rect 9655 51113 9689 51147
rect 9991 51113 10025 51147
rect 10327 51113 10361 51147
rect 10663 51113 10697 51147
rect 10999 51113 11033 51147
rect 11335 51113 11369 51147
rect 11671 51113 11705 51147
rect 12007 51113 12041 51147
rect 12343 51113 12377 51147
rect 12679 51113 12713 51147
rect 13015 51113 13049 51147
rect 13351 51113 13385 51147
rect 13687 51113 13721 51147
rect 14023 51113 14057 51147
rect 14359 51113 14393 51147
rect 14695 51113 14729 51147
rect 15031 51113 15065 51147
rect 15367 51113 15401 51147
rect 15703 51113 15737 51147
rect 16039 51113 16073 51147
rect 16375 51113 16409 51147
rect 16711 51113 16745 51147
rect 17047 51113 17081 51147
rect 17383 51113 17417 51147
rect 17719 51113 17753 51147
rect 18055 51113 18089 51147
rect 18391 51113 18425 51147
rect 18727 51113 18761 51147
rect 19063 51113 19097 51147
rect 19399 51113 19433 51147
rect 19735 51113 19769 51147
rect 20071 51113 20105 51147
rect 20407 51113 20441 51147
rect 20743 51113 20777 51147
rect 21079 51113 21113 51147
rect 21415 51113 21449 51147
rect 21751 51113 21785 51147
rect 22087 51113 22121 51147
rect 22423 51113 22457 51147
rect 22759 51113 22793 51147
rect 23095 51113 23129 51147
rect 23431 51113 23465 51147
rect 23767 51113 23801 51147
rect 24103 51113 24137 51147
rect 24439 51113 24473 51147
rect 24775 51113 24809 51147
rect 25111 51113 25145 51147
rect 25447 51113 25481 51147
rect 25783 51113 25817 51147
rect 26119 51113 26153 51147
rect 26455 51113 26489 51147
rect 26791 51113 26825 51147
rect 27127 51113 27161 51147
rect 27463 51113 27497 51147
rect 27799 51113 27833 51147
rect 28135 51113 28169 51147
rect 28471 51113 28505 51147
rect 28807 51113 28841 51147
rect 29143 51113 29177 51147
rect 29479 51113 29513 51147
rect 29815 51113 29849 51147
rect 30151 51113 30185 51147
rect 30487 51113 30521 51147
rect 30823 51113 30857 51147
rect 31159 51113 31193 51147
rect 31495 51113 31529 51147
rect 31831 51113 31865 51147
rect 32167 51113 32201 51147
rect 32503 51113 32537 51147
rect 32839 51113 32873 51147
rect 33175 51113 33209 51147
rect 33511 51113 33545 51147
rect 33847 51113 33881 51147
rect 34183 51113 34217 51147
rect 34519 51113 34553 51147
rect 34855 51113 34889 51147
rect 35191 51113 35225 51147
rect 35527 51113 35561 51147
rect 35863 51113 35897 51147
rect 36199 51113 36233 51147
rect 36535 51113 36569 51147
rect 36871 51113 36905 51147
rect 37207 51113 37241 51147
rect 37543 51113 37577 51147
rect 37879 51113 37913 51147
rect 38215 51113 38249 51147
rect 38551 51113 38585 51147
rect 38887 51113 38921 51147
rect 39223 51113 39257 51147
rect 39559 51113 39593 51147
rect 39895 51113 39929 51147
rect 40231 51113 40265 51147
rect 40567 51113 40601 51147
rect 40903 51113 40937 51147
rect 41239 51113 41273 51147
rect 41575 51113 41609 51147
rect 41911 51113 41945 51147
rect 42247 51113 42281 51147
rect 42583 51113 42617 51147
rect 42919 51113 42953 51147
rect 43255 51113 43289 51147
rect 43591 51113 43625 51147
rect 43927 51113 43961 51147
rect 44263 51113 44297 51147
rect 44599 51113 44633 51147
rect 44935 51113 44969 51147
rect 45271 51113 45305 51147
rect 45607 51113 45641 51147
rect 45943 51113 45977 51147
rect 46279 51113 46313 51147
rect 46615 51113 46649 51147
rect 46951 51113 46985 51147
rect 47287 51113 47321 51147
rect 47623 51113 47657 51147
rect 47959 51113 47993 51147
rect 48295 51113 48329 51147
rect 48631 51113 48665 51147
rect 48967 51113 49001 51147
rect 49303 51113 49337 51147
rect 49639 51113 49673 51147
rect 49975 51113 50009 51147
rect 50311 51113 50345 51147
rect 50647 51113 50681 51147
rect 50983 51113 51017 51147
rect 51319 51113 51353 51147
rect 51655 51113 51689 51147
rect 51991 51113 52025 51147
rect 52327 51113 52361 51147
rect 52663 51113 52697 51147
rect 52999 51113 53033 51147
rect 53335 51113 53369 51147
rect 53671 51113 53705 51147
rect 54007 51113 54041 51147
rect 54343 51113 54377 51147
rect 54679 51113 54713 51147
rect 55015 51113 55049 51147
rect 55351 51113 55385 51147
rect 55687 51113 55721 51147
rect 56023 51113 56057 51147
rect 56359 51113 56393 51147
rect 56695 51113 56729 51147
rect 57031 51113 57065 51147
rect 57367 51113 57401 51147
rect 57703 51113 57737 51147
rect 58039 51113 58073 51147
rect 58375 51113 58409 51147
rect 58711 51113 58745 51147
rect 59047 51113 59081 51147
rect 59383 51113 59417 51147
rect 59719 51113 59753 51147
rect 60055 51113 60089 51147
rect 60391 51113 60425 51147
rect 60727 51113 60761 51147
rect 61063 51113 61097 51147
rect 61399 51113 61433 51147
rect 61735 51113 61769 51147
rect 62071 51113 62105 51147
rect 62407 51113 62441 51147
rect 62743 51113 62777 51147
rect 63079 51113 63113 51147
rect 63415 51113 63449 51147
rect 63751 51113 63785 51147
rect 64087 51113 64121 51147
rect 64423 51113 64457 51147
rect 64759 51113 64793 51147
rect 65095 51113 65129 51147
rect 65431 51113 65465 51147
rect 65767 51113 65801 51147
rect 1591 50647 1625 50681
rect 66195 50647 66229 50681
rect 1591 50311 1625 50345
rect 66195 50311 66229 50345
rect 1591 49975 1625 50009
rect 66195 49975 66229 50009
rect 1591 49639 1625 49673
rect 66195 49639 66229 49673
rect 1591 49303 1625 49337
rect 66195 49303 66229 49337
rect 1591 48967 1625 49001
rect 66195 48967 66229 49001
rect 1591 48631 1625 48665
rect 66195 48631 66229 48665
rect 1591 48295 1625 48329
rect 66195 48295 66229 48329
rect 1591 47959 1625 47993
rect 66195 47959 66229 47993
rect 1591 47623 1625 47657
rect 66195 47623 66229 47657
rect 1591 47287 1625 47321
rect 66195 47287 66229 47321
rect 1591 46951 1625 46985
rect 66195 46951 66229 46985
rect 1591 46615 1625 46649
rect 66195 46615 66229 46649
rect 1591 46279 1625 46313
rect 66195 46279 66229 46313
rect 1591 45943 1625 45977
rect 66195 45943 66229 45977
rect 1591 45607 1625 45641
rect 66195 45607 66229 45641
rect 1591 45271 1625 45305
rect 66195 45271 66229 45305
rect 1591 44935 1625 44969
rect 66195 44935 66229 44969
rect 1591 44599 1625 44633
rect 66195 44599 66229 44633
rect 1591 44263 1625 44297
rect 66195 44263 66229 44297
rect 1591 43927 1625 43961
rect 66195 43927 66229 43961
rect 1591 43591 1625 43625
rect 66195 43591 66229 43625
rect 1591 43255 1625 43289
rect 66195 43255 66229 43289
rect 1591 42919 1625 42953
rect 66195 42919 66229 42953
rect 1591 42583 1625 42617
rect 66195 42583 66229 42617
rect 1591 42247 1625 42281
rect 66195 42247 66229 42281
rect 1591 41911 1625 41945
rect 66195 41911 66229 41945
rect 1591 41575 1625 41609
rect 66195 41575 66229 41609
rect 1591 41239 1625 41273
rect 66195 41239 66229 41273
rect 1591 40903 1625 40937
rect 66195 40903 66229 40937
rect 1591 40567 1625 40601
rect 66195 40567 66229 40601
rect 1591 40231 1625 40265
rect 66195 40231 66229 40265
rect 1591 39895 1625 39929
rect 66195 39895 66229 39929
rect 1591 39559 1625 39593
rect 66195 39559 66229 39593
rect 1591 39223 1625 39257
rect 66195 39223 66229 39257
rect 1591 38887 1625 38921
rect 66195 38887 66229 38921
rect 1591 38551 1625 38585
rect 66195 38551 66229 38585
rect 1591 38215 1625 38249
rect 66195 38215 66229 38249
rect 1591 37879 1625 37913
rect 66195 37879 66229 37913
rect 1591 37543 1625 37577
rect 66195 37543 66229 37577
rect 1591 37207 1625 37241
rect 66195 37207 66229 37241
rect 1591 36871 1625 36905
rect 66195 36871 66229 36905
rect 1591 36535 1625 36569
rect 66195 36535 66229 36569
rect 1591 36199 1625 36233
rect 66195 36199 66229 36233
rect 1591 35863 1625 35897
rect 66195 35863 66229 35897
rect 1591 35527 1625 35561
rect 66195 35527 66229 35561
rect 1591 35191 1625 35225
rect 66195 35191 66229 35225
rect 1591 34855 1625 34889
rect 66195 34855 66229 34889
rect 1591 34519 1625 34553
rect 66195 34519 66229 34553
rect 1591 34183 1625 34217
rect 66195 34183 66229 34217
rect 1591 33847 1625 33881
rect 66195 33847 66229 33881
rect 1591 33511 1625 33545
rect 66195 33511 66229 33545
rect 1591 33175 1625 33209
rect 66195 33175 66229 33209
rect 1591 32839 1625 32873
rect 66195 32839 66229 32873
rect 1591 32503 1625 32537
rect 66195 32503 66229 32537
rect 1591 32167 1625 32201
rect 66195 32167 66229 32201
rect 1591 31831 1625 31865
rect 66195 31831 66229 31865
rect 1591 31495 1625 31529
rect 66195 31495 66229 31529
rect 1591 31159 1625 31193
rect 66195 31159 66229 31193
rect 1591 30823 1625 30857
rect 66195 30823 66229 30857
rect 1591 30487 1625 30521
rect 66195 30487 66229 30521
rect 1591 30151 1625 30185
rect 66195 30151 66229 30185
rect 1591 29815 1625 29849
rect 66195 29815 66229 29849
rect 1591 29479 1625 29513
rect 66195 29479 66229 29513
rect 1591 29143 1625 29177
rect 66195 29143 66229 29177
rect 1591 28807 1625 28841
rect 66195 28807 66229 28841
rect 1591 28471 1625 28505
rect 66195 28471 66229 28505
rect 1591 28135 1625 28169
rect 66195 28135 66229 28169
rect 1591 27799 1625 27833
rect 66195 27799 66229 27833
rect 1591 27463 1625 27497
rect 66195 27463 66229 27497
rect 1591 27127 1625 27161
rect 66195 27127 66229 27161
rect 1591 26791 1625 26825
rect 66195 26791 66229 26825
rect 1591 26455 1625 26489
rect 66195 26455 66229 26489
rect 1591 26119 1625 26153
rect 66195 26119 66229 26153
rect 1591 25783 1625 25817
rect 66195 25783 66229 25817
rect 1591 25447 1625 25481
rect 66195 25447 66229 25481
rect 1591 25111 1625 25145
rect 66195 25111 66229 25145
rect 1591 24775 1625 24809
rect 66195 24775 66229 24809
rect 1591 24439 1625 24473
rect 66195 24439 66229 24473
rect 1591 24103 1625 24137
rect 66195 24103 66229 24137
rect 1591 23767 1625 23801
rect 66195 23767 66229 23801
rect 1591 23431 1625 23465
rect 66195 23431 66229 23465
rect 1591 23095 1625 23129
rect 66195 23095 66229 23129
rect 1591 22759 1625 22793
rect 66195 22759 66229 22793
rect 1591 22423 1625 22457
rect 66195 22423 66229 22457
rect 1591 22087 1625 22121
rect 66195 22087 66229 22121
rect 1591 21751 1625 21785
rect 66195 21751 66229 21785
rect 1591 21415 1625 21449
rect 66195 21415 66229 21449
rect 1591 21079 1625 21113
rect 66195 21079 66229 21113
rect 1591 20743 1625 20777
rect 66195 20743 66229 20777
rect 1591 20407 1625 20441
rect 66195 20407 66229 20441
rect 1591 20071 1625 20105
rect 66195 20071 66229 20105
rect 1591 19735 1625 19769
rect 66195 19735 66229 19769
rect 1591 19399 1625 19433
rect 66195 19399 66229 19433
rect 1591 19063 1625 19097
rect 66195 19063 66229 19097
rect 1591 18727 1625 18761
rect 66195 18727 66229 18761
rect 1591 18391 1625 18425
rect 66195 18391 66229 18425
rect 1591 18055 1625 18089
rect 66195 18055 66229 18089
rect 1591 17719 1625 17753
rect 66195 17719 66229 17753
rect 1591 17383 1625 17417
rect 66195 17383 66229 17417
rect 1591 17047 1625 17081
rect 66195 17047 66229 17081
rect 1591 16711 1625 16745
rect 66195 16711 66229 16745
rect 1591 16375 1625 16409
rect 66195 16375 66229 16409
rect 1591 16039 1625 16073
rect 66195 16039 66229 16073
rect 1591 15703 1625 15737
rect 66195 15703 66229 15737
rect 1591 15367 1625 15401
rect 66195 15367 66229 15401
rect 1591 15031 1625 15065
rect 66195 15031 66229 15065
rect 1591 14695 1625 14729
rect 66195 14695 66229 14729
rect 1591 14359 1625 14393
rect 66195 14359 66229 14393
rect 1591 14023 1625 14057
rect 66195 14023 66229 14057
rect 1591 13687 1625 13721
rect 66195 13687 66229 13721
rect 1591 13351 1625 13385
rect 66195 13351 66229 13385
rect 1591 13015 1625 13049
rect 66195 13015 66229 13049
rect 1591 12679 1625 12713
rect 66195 12679 66229 12713
rect 1591 12343 1625 12377
rect 66195 12343 66229 12377
rect 1591 12007 1625 12041
rect 66195 12007 66229 12041
rect 1591 11671 1625 11705
rect 66195 11671 66229 11705
rect 1591 11335 1625 11369
rect 66195 11335 66229 11369
rect 1591 10999 1625 11033
rect 66195 10999 66229 11033
rect 1591 10663 1625 10697
rect 66195 10663 66229 10697
rect 1591 10327 1625 10361
rect 66195 10327 66229 10361
rect 1591 9991 1625 10025
rect 66195 9991 66229 10025
rect 1591 9655 1625 9689
rect 66195 9655 66229 9689
rect 1591 9319 1625 9353
rect 66195 9319 66229 9353
rect 1591 8983 1625 9017
rect 66195 8983 66229 9017
rect 1591 8647 1625 8681
rect 66195 8647 66229 8681
rect 1591 8311 1625 8345
rect 66195 8311 66229 8345
rect 1591 7975 1625 8009
rect 66195 7975 66229 8009
rect 1591 7639 1625 7673
rect 66195 7639 66229 7673
rect 1591 7303 1625 7337
rect 66195 7303 66229 7337
rect 1591 6967 1625 7001
rect 66195 6967 66229 7001
rect 1591 6631 1625 6665
rect 66195 6631 66229 6665
rect 1591 6295 1625 6329
rect 66195 6295 66229 6329
rect 1591 5959 1625 5993
rect 66195 5959 66229 5993
rect 1591 5623 1625 5657
rect 66195 5623 66229 5657
rect 1591 5287 1625 5321
rect 66195 5287 66229 5321
rect 1591 4951 1625 4985
rect 66195 4951 66229 4985
rect 1591 4615 1625 4649
rect 66195 4615 66229 4649
rect 1591 4279 1625 4313
rect 66195 4279 66229 4313
rect 1591 3943 1625 3977
rect 66195 3943 66229 3977
rect 1591 3607 1625 3641
rect 66195 3607 66229 3641
rect 1591 3271 1625 3305
rect 66195 3271 66229 3305
rect 1591 2935 1625 2969
rect 66195 2935 66229 2969
rect 1591 2599 1625 2633
rect 66195 2599 66229 2633
rect 1591 2263 1625 2297
rect 66195 2263 66229 2297
rect 1591 1927 1625 1961
rect 66195 1927 66229 1961
rect 1927 1591 1961 1625
rect 2263 1591 2297 1625
rect 2599 1591 2633 1625
rect 2935 1591 2969 1625
rect 3271 1591 3305 1625
rect 3607 1591 3641 1625
rect 3943 1591 3977 1625
rect 4279 1591 4313 1625
rect 4615 1591 4649 1625
rect 4951 1591 4985 1625
rect 5287 1591 5321 1625
rect 5623 1591 5657 1625
rect 5959 1591 5993 1625
rect 6295 1591 6329 1625
rect 6631 1591 6665 1625
rect 6967 1591 7001 1625
rect 7303 1591 7337 1625
rect 7639 1591 7673 1625
rect 7975 1591 8009 1625
rect 8311 1591 8345 1625
rect 8647 1591 8681 1625
rect 8983 1591 9017 1625
rect 9319 1591 9353 1625
rect 9655 1591 9689 1625
rect 9991 1591 10025 1625
rect 10327 1591 10361 1625
rect 10663 1591 10697 1625
rect 10999 1591 11033 1625
rect 11335 1591 11369 1625
rect 11671 1591 11705 1625
rect 12007 1591 12041 1625
rect 12343 1591 12377 1625
rect 12679 1591 12713 1625
rect 13015 1591 13049 1625
rect 13351 1591 13385 1625
rect 13687 1591 13721 1625
rect 14023 1591 14057 1625
rect 14359 1591 14393 1625
rect 14695 1591 14729 1625
rect 15031 1591 15065 1625
rect 15367 1591 15401 1625
rect 15703 1591 15737 1625
rect 16039 1591 16073 1625
rect 16375 1591 16409 1625
rect 16711 1591 16745 1625
rect 17047 1591 17081 1625
rect 17383 1591 17417 1625
rect 17719 1591 17753 1625
rect 18055 1591 18089 1625
rect 18391 1591 18425 1625
rect 18727 1591 18761 1625
rect 19063 1591 19097 1625
rect 19399 1591 19433 1625
rect 19735 1591 19769 1625
rect 20071 1591 20105 1625
rect 20407 1591 20441 1625
rect 20743 1591 20777 1625
rect 21079 1591 21113 1625
rect 21415 1591 21449 1625
rect 21751 1591 21785 1625
rect 22087 1591 22121 1625
rect 22423 1591 22457 1625
rect 22759 1591 22793 1625
rect 23095 1591 23129 1625
rect 23431 1591 23465 1625
rect 23767 1591 23801 1625
rect 24103 1591 24137 1625
rect 24439 1591 24473 1625
rect 24775 1591 24809 1625
rect 25111 1591 25145 1625
rect 25447 1591 25481 1625
rect 25783 1591 25817 1625
rect 26119 1591 26153 1625
rect 26455 1591 26489 1625
rect 26791 1591 26825 1625
rect 27127 1591 27161 1625
rect 27463 1591 27497 1625
rect 27799 1591 27833 1625
rect 28135 1591 28169 1625
rect 28471 1591 28505 1625
rect 28807 1591 28841 1625
rect 29143 1591 29177 1625
rect 29479 1591 29513 1625
rect 29815 1591 29849 1625
rect 30151 1591 30185 1625
rect 30487 1591 30521 1625
rect 30823 1591 30857 1625
rect 31159 1591 31193 1625
rect 31495 1591 31529 1625
rect 31831 1591 31865 1625
rect 32167 1591 32201 1625
rect 32503 1591 32537 1625
rect 32839 1591 32873 1625
rect 33175 1591 33209 1625
rect 33511 1591 33545 1625
rect 33847 1591 33881 1625
rect 34183 1591 34217 1625
rect 34519 1591 34553 1625
rect 34855 1591 34889 1625
rect 35191 1591 35225 1625
rect 35527 1591 35561 1625
rect 35863 1591 35897 1625
rect 36199 1591 36233 1625
rect 36535 1591 36569 1625
rect 36871 1591 36905 1625
rect 37207 1591 37241 1625
rect 37543 1591 37577 1625
rect 37879 1591 37913 1625
rect 38215 1591 38249 1625
rect 38551 1591 38585 1625
rect 38887 1591 38921 1625
rect 39223 1591 39257 1625
rect 39559 1591 39593 1625
rect 39895 1591 39929 1625
rect 40231 1591 40265 1625
rect 40567 1591 40601 1625
rect 40903 1591 40937 1625
rect 41239 1591 41273 1625
rect 41575 1591 41609 1625
rect 41911 1591 41945 1625
rect 42247 1591 42281 1625
rect 42583 1591 42617 1625
rect 42919 1591 42953 1625
rect 43255 1591 43289 1625
rect 43591 1591 43625 1625
rect 43927 1591 43961 1625
rect 44263 1591 44297 1625
rect 44599 1591 44633 1625
rect 44935 1591 44969 1625
rect 45271 1591 45305 1625
rect 45607 1591 45641 1625
rect 45943 1591 45977 1625
rect 46279 1591 46313 1625
rect 46615 1591 46649 1625
rect 46951 1591 46985 1625
rect 47287 1591 47321 1625
rect 47623 1591 47657 1625
rect 47959 1591 47993 1625
rect 48295 1591 48329 1625
rect 48631 1591 48665 1625
rect 48967 1591 49001 1625
rect 49303 1591 49337 1625
rect 49639 1591 49673 1625
rect 49975 1591 50009 1625
rect 50311 1591 50345 1625
rect 50647 1591 50681 1625
rect 50983 1591 51017 1625
rect 51319 1591 51353 1625
rect 51655 1591 51689 1625
rect 51991 1591 52025 1625
rect 52327 1591 52361 1625
rect 52663 1591 52697 1625
rect 52999 1591 53033 1625
rect 53335 1591 53369 1625
rect 53671 1591 53705 1625
rect 54007 1591 54041 1625
rect 54343 1591 54377 1625
rect 54679 1591 54713 1625
rect 55015 1591 55049 1625
rect 55351 1591 55385 1625
rect 55687 1591 55721 1625
rect 56023 1591 56057 1625
rect 56359 1591 56393 1625
rect 56695 1591 56729 1625
rect 57031 1591 57065 1625
rect 57367 1591 57401 1625
rect 57703 1591 57737 1625
rect 58039 1591 58073 1625
rect 58375 1591 58409 1625
rect 58711 1591 58745 1625
rect 59047 1591 59081 1625
rect 59383 1591 59417 1625
rect 59719 1591 59753 1625
rect 60055 1591 60089 1625
rect 60391 1591 60425 1625
rect 60727 1591 60761 1625
rect 61063 1591 61097 1625
rect 61399 1591 61433 1625
rect 61735 1591 61769 1625
rect 62071 1591 62105 1625
rect 62407 1591 62441 1625
rect 62743 1591 62777 1625
rect 63079 1591 63113 1625
rect 63415 1591 63449 1625
rect 63751 1591 63785 1625
rect 64087 1591 64121 1625
rect 64423 1591 64457 1625
rect 64759 1591 64793 1625
rect 65095 1591 65129 1625
rect 65431 1591 65465 1625
rect 65767 1591 65801 1625
<< metal1 >>
rect 1496 51156 66324 51242
rect 1496 51104 1918 51156
rect 1970 51147 3598 51156
rect 3650 51147 5278 51156
rect 5330 51147 6958 51156
rect 7010 51147 8638 51156
rect 8690 51147 10318 51156
rect 10370 51147 11998 51156
rect 12050 51147 13678 51156
rect 13730 51147 15358 51156
rect 15410 51147 17038 51156
rect 17090 51147 18718 51156
rect 18770 51147 20398 51156
rect 20450 51147 22078 51156
rect 22130 51147 23758 51156
rect 23810 51147 25438 51156
rect 25490 51147 27118 51156
rect 27170 51147 28798 51156
rect 28850 51147 30478 51156
rect 30530 51147 32158 51156
rect 32210 51147 33838 51156
rect 33890 51147 35518 51156
rect 35570 51147 37198 51156
rect 37250 51147 38878 51156
rect 38930 51147 40558 51156
rect 40610 51147 42238 51156
rect 42290 51147 43918 51156
rect 43970 51147 45598 51156
rect 45650 51147 47278 51156
rect 47330 51147 48958 51156
rect 49010 51147 50638 51156
rect 50690 51147 52318 51156
rect 52370 51147 53998 51156
rect 54050 51147 55678 51156
rect 55730 51147 57358 51156
rect 57410 51147 59038 51156
rect 59090 51147 60718 51156
rect 60770 51147 62398 51156
rect 62450 51147 64078 51156
rect 64130 51147 65758 51156
rect 1970 51113 2263 51147
rect 2297 51113 2599 51147
rect 2633 51113 2935 51147
rect 2969 51113 3271 51147
rect 3305 51113 3598 51147
rect 3650 51113 3943 51147
rect 3977 51113 4279 51147
rect 4313 51113 4615 51147
rect 4649 51113 4951 51147
rect 4985 51113 5278 51147
rect 5330 51113 5623 51147
rect 5657 51113 5959 51147
rect 5993 51113 6295 51147
rect 6329 51113 6631 51147
rect 6665 51113 6958 51147
rect 7010 51113 7303 51147
rect 7337 51113 7639 51147
rect 7673 51113 7975 51147
rect 8009 51113 8311 51147
rect 8345 51113 8638 51147
rect 8690 51113 8983 51147
rect 9017 51113 9319 51147
rect 9353 51113 9655 51147
rect 9689 51113 9991 51147
rect 10025 51113 10318 51147
rect 10370 51113 10663 51147
rect 10697 51113 10999 51147
rect 11033 51113 11335 51147
rect 11369 51113 11671 51147
rect 11705 51113 11998 51147
rect 12050 51113 12343 51147
rect 12377 51113 12679 51147
rect 12713 51113 13015 51147
rect 13049 51113 13351 51147
rect 13385 51113 13678 51147
rect 13730 51113 14023 51147
rect 14057 51113 14359 51147
rect 14393 51113 14695 51147
rect 14729 51113 15031 51147
rect 15065 51113 15358 51147
rect 15410 51113 15703 51147
rect 15737 51113 16039 51147
rect 16073 51113 16375 51147
rect 16409 51113 16711 51147
rect 16745 51113 17038 51147
rect 17090 51113 17383 51147
rect 17417 51113 17719 51147
rect 17753 51113 18055 51147
rect 18089 51113 18391 51147
rect 18425 51113 18718 51147
rect 18770 51113 19063 51147
rect 19097 51113 19399 51147
rect 19433 51113 19735 51147
rect 19769 51113 20071 51147
rect 20105 51113 20398 51147
rect 20450 51113 20743 51147
rect 20777 51113 21079 51147
rect 21113 51113 21415 51147
rect 21449 51113 21751 51147
rect 21785 51113 22078 51147
rect 22130 51113 22423 51147
rect 22457 51113 22759 51147
rect 22793 51113 23095 51147
rect 23129 51113 23431 51147
rect 23465 51113 23758 51147
rect 23810 51113 24103 51147
rect 24137 51113 24439 51147
rect 24473 51113 24775 51147
rect 24809 51113 25111 51147
rect 25145 51113 25438 51147
rect 25490 51113 25783 51147
rect 25817 51113 26119 51147
rect 26153 51113 26455 51147
rect 26489 51113 26791 51147
rect 26825 51113 27118 51147
rect 27170 51113 27463 51147
rect 27497 51113 27799 51147
rect 27833 51113 28135 51147
rect 28169 51113 28471 51147
rect 28505 51113 28798 51147
rect 28850 51113 29143 51147
rect 29177 51113 29479 51147
rect 29513 51113 29815 51147
rect 29849 51113 30151 51147
rect 30185 51113 30478 51147
rect 30530 51113 30823 51147
rect 30857 51113 31159 51147
rect 31193 51113 31495 51147
rect 31529 51113 31831 51147
rect 31865 51113 32158 51147
rect 32210 51113 32503 51147
rect 32537 51113 32839 51147
rect 32873 51113 33175 51147
rect 33209 51113 33511 51147
rect 33545 51113 33838 51147
rect 33890 51113 34183 51147
rect 34217 51113 34519 51147
rect 34553 51113 34855 51147
rect 34889 51113 35191 51147
rect 35225 51113 35518 51147
rect 35570 51113 35863 51147
rect 35897 51113 36199 51147
rect 36233 51113 36535 51147
rect 36569 51113 36871 51147
rect 36905 51113 37198 51147
rect 37250 51113 37543 51147
rect 37577 51113 37879 51147
rect 37913 51113 38215 51147
rect 38249 51113 38551 51147
rect 38585 51113 38878 51147
rect 38930 51113 39223 51147
rect 39257 51113 39559 51147
rect 39593 51113 39895 51147
rect 39929 51113 40231 51147
rect 40265 51113 40558 51147
rect 40610 51113 40903 51147
rect 40937 51113 41239 51147
rect 41273 51113 41575 51147
rect 41609 51113 41911 51147
rect 41945 51113 42238 51147
rect 42290 51113 42583 51147
rect 42617 51113 42919 51147
rect 42953 51113 43255 51147
rect 43289 51113 43591 51147
rect 43625 51113 43918 51147
rect 43970 51113 44263 51147
rect 44297 51113 44599 51147
rect 44633 51113 44935 51147
rect 44969 51113 45271 51147
rect 45305 51113 45598 51147
rect 45650 51113 45943 51147
rect 45977 51113 46279 51147
rect 46313 51113 46615 51147
rect 46649 51113 46951 51147
rect 46985 51113 47278 51147
rect 47330 51113 47623 51147
rect 47657 51113 47959 51147
rect 47993 51113 48295 51147
rect 48329 51113 48631 51147
rect 48665 51113 48958 51147
rect 49010 51113 49303 51147
rect 49337 51113 49639 51147
rect 49673 51113 49975 51147
rect 50009 51113 50311 51147
rect 50345 51113 50638 51147
rect 50690 51113 50983 51147
rect 51017 51113 51319 51147
rect 51353 51113 51655 51147
rect 51689 51113 51991 51147
rect 52025 51113 52318 51147
rect 52370 51113 52663 51147
rect 52697 51113 52999 51147
rect 53033 51113 53335 51147
rect 53369 51113 53671 51147
rect 53705 51113 53998 51147
rect 54050 51113 54343 51147
rect 54377 51113 54679 51147
rect 54713 51113 55015 51147
rect 55049 51113 55351 51147
rect 55385 51113 55678 51147
rect 55730 51113 56023 51147
rect 56057 51113 56359 51147
rect 56393 51113 56695 51147
rect 56729 51113 57031 51147
rect 57065 51113 57358 51147
rect 57410 51113 57703 51147
rect 57737 51113 58039 51147
rect 58073 51113 58375 51147
rect 58409 51113 58711 51147
rect 58745 51113 59038 51147
rect 59090 51113 59383 51147
rect 59417 51113 59719 51147
rect 59753 51113 60055 51147
rect 60089 51113 60391 51147
rect 60425 51113 60718 51147
rect 60770 51113 61063 51147
rect 61097 51113 61399 51147
rect 61433 51113 61735 51147
rect 61769 51113 62071 51147
rect 62105 51113 62398 51147
rect 62450 51113 62743 51147
rect 62777 51113 63079 51147
rect 63113 51113 63415 51147
rect 63449 51113 63751 51147
rect 63785 51113 64078 51147
rect 64130 51113 64423 51147
rect 64457 51113 64759 51147
rect 64793 51113 65095 51147
rect 65129 51113 65431 51147
rect 65465 51113 65758 51147
rect 1970 51104 3598 51113
rect 3650 51104 5278 51113
rect 5330 51104 6958 51113
rect 7010 51104 8638 51113
rect 8690 51104 10318 51113
rect 10370 51104 11998 51113
rect 12050 51104 13678 51113
rect 13730 51104 15358 51113
rect 15410 51104 17038 51113
rect 17090 51104 18718 51113
rect 18770 51104 20398 51113
rect 20450 51104 22078 51113
rect 22130 51104 23758 51113
rect 23810 51104 25438 51113
rect 25490 51104 27118 51113
rect 27170 51104 28798 51113
rect 28850 51104 30478 51113
rect 30530 51104 32158 51113
rect 32210 51104 33838 51113
rect 33890 51104 35518 51113
rect 35570 51104 37198 51113
rect 37250 51104 38878 51113
rect 38930 51104 40558 51113
rect 40610 51104 42238 51113
rect 42290 51104 43918 51113
rect 43970 51104 45598 51113
rect 45650 51104 47278 51113
rect 47330 51104 48958 51113
rect 49010 51104 50638 51113
rect 50690 51104 52318 51113
rect 52370 51104 53998 51113
rect 54050 51104 55678 51113
rect 55730 51104 57358 51113
rect 57410 51104 59038 51113
rect 59090 51104 60718 51113
rect 60770 51104 62398 51113
rect 62450 51104 64078 51113
rect 64130 51104 65758 51113
rect 65810 51104 66324 51156
rect 1496 51018 66324 51104
rect 1576 50638 1582 50690
rect 1634 50638 1640 50690
rect 66180 50638 66186 50690
rect 66238 50638 66244 50690
rect 1576 50302 1582 50354
rect 1634 50302 1640 50354
rect 66180 50302 66186 50354
rect 66238 50302 66244 50354
rect 1576 49966 1582 50018
rect 1634 49966 1640 50018
rect 66180 49966 66186 50018
rect 66238 49966 66244 50018
rect 1576 49630 1582 49682
rect 1634 49630 1640 49682
rect 66180 49630 66186 49682
rect 66238 49630 66244 49682
rect 1576 49294 1582 49346
rect 1634 49294 1640 49346
rect 66180 49294 66186 49346
rect 66238 49294 66244 49346
rect 1576 48958 1582 49010
rect 1634 48958 1640 49010
rect 66180 48958 66186 49010
rect 66238 48958 66244 49010
rect 1576 48622 1582 48674
rect 1634 48622 1640 48674
rect 66180 48622 66186 48674
rect 66238 48622 66244 48674
rect 1576 48286 1582 48338
rect 1634 48286 1640 48338
rect 66180 48286 66186 48338
rect 66238 48286 66244 48338
rect 1576 47950 1582 48002
rect 1634 47950 1640 48002
rect 66180 47950 66186 48002
rect 66238 47950 66244 48002
rect 1576 47614 1582 47666
rect 1634 47614 1640 47666
rect 66180 47614 66186 47666
rect 66238 47614 66244 47666
rect 1576 47278 1582 47330
rect 1634 47278 1640 47330
rect 66180 47278 66186 47330
rect 66238 47278 66244 47330
rect 1576 46942 1582 46994
rect 1634 46942 1640 46994
rect 66180 46942 66186 46994
rect 66238 46942 66244 46994
rect 23979 46835 23985 46887
rect 24037 46835 24043 46887
rect 26475 46835 26481 46887
rect 26533 46835 26539 46887
rect 28971 46835 28977 46887
rect 29029 46835 29035 46887
rect 31467 46835 31473 46887
rect 31525 46835 31531 46887
rect 33963 46835 33969 46887
rect 34021 46835 34027 46887
rect 36459 46835 36465 46887
rect 36517 46835 36523 46887
rect 38955 46835 38961 46887
rect 39013 46835 39019 46887
rect 41451 46835 41457 46887
rect 41509 46835 41515 46887
rect 1576 46606 1582 46658
rect 1634 46606 1640 46658
rect 66180 46606 66186 46658
rect 66238 46606 66244 46658
rect 1576 46270 1582 46322
rect 1634 46270 1640 46322
rect 66180 46270 66186 46322
rect 66238 46270 66244 46322
rect 1576 45934 1582 45986
rect 1634 45934 1640 45986
rect 66180 45934 66186 45986
rect 66238 45934 66244 45986
rect 1576 45598 1582 45650
rect 1634 45598 1640 45650
rect 66180 45598 66186 45650
rect 66238 45598 66244 45650
rect 1576 45262 1582 45314
rect 1634 45262 1640 45314
rect 66180 45262 66186 45314
rect 66238 45262 66244 45314
rect 1576 44926 1582 44978
rect 1634 44926 1640 44978
rect 66180 44926 66186 44978
rect 66238 44926 66244 44978
rect 1576 44590 1582 44642
rect 1634 44590 1640 44642
rect 66180 44590 66186 44642
rect 66238 44590 66244 44642
rect 1576 44254 1582 44306
rect 1634 44254 1640 44306
rect 66180 44254 66186 44306
rect 66238 44254 66244 44306
rect 1576 43918 1582 43970
rect 1634 43918 1640 43970
rect 66180 43918 66186 43970
rect 66238 43918 66244 43970
rect 1576 43582 1582 43634
rect 1634 43582 1640 43634
rect 66180 43582 66186 43634
rect 66238 43582 66244 43634
rect 1576 43246 1582 43298
rect 1634 43246 1640 43298
rect 66180 43246 66186 43298
rect 66238 43246 66244 43298
rect 1576 42910 1582 42962
rect 1634 42910 1640 42962
rect 66180 42910 66186 42962
rect 66238 42910 66244 42962
rect 1576 42574 1582 42626
rect 1634 42574 1640 42626
rect 66180 42574 66186 42626
rect 66238 42574 66244 42626
rect 1576 42238 1582 42290
rect 1634 42238 1640 42290
rect 66180 42238 66186 42290
rect 66238 42238 66244 42290
rect 1576 41902 1582 41954
rect 1634 41902 1640 41954
rect 66180 41902 66186 41954
rect 66238 41902 66244 41954
rect 1576 41566 1582 41618
rect 1634 41566 1640 41618
rect 66180 41566 66186 41618
rect 66238 41566 66244 41618
rect 1576 41230 1582 41282
rect 1634 41230 1640 41282
rect 66180 41230 66186 41282
rect 66238 41230 66244 41282
rect 1576 40894 1582 40946
rect 1634 40894 1640 40946
rect 66180 40894 66186 40946
rect 66238 40894 66244 40946
rect 1576 40558 1582 40610
rect 1634 40558 1640 40610
rect 66180 40558 66186 40610
rect 66238 40558 66244 40610
rect 1576 40222 1582 40274
rect 1634 40222 1640 40274
rect 66180 40222 66186 40274
rect 66238 40222 66244 40274
rect 46765 40100 46771 40152
rect 46823 40100 46829 40152
rect 48656 40087 48662 40139
rect 48714 40087 48720 40139
rect 1576 39886 1582 39938
rect 1634 39886 1640 39938
rect 66180 39886 66186 39938
rect 66238 39886 66244 39938
rect 1576 39550 1582 39602
rect 1634 39550 1640 39602
rect 66180 39550 66186 39602
rect 66238 39550 66244 39602
rect 1576 39214 1582 39266
rect 1634 39214 1640 39266
rect 66180 39214 66186 39266
rect 66238 39214 66244 39266
rect 1576 38878 1582 38930
rect 1634 38878 1640 38930
rect 66180 38878 66186 38930
rect 66238 38878 66244 38930
rect 1576 38542 1582 38594
rect 1634 38542 1640 38594
rect 66180 38542 66186 38594
rect 66238 38542 66244 38594
rect 1576 38206 1582 38258
rect 1634 38206 1640 38258
rect 66180 38206 66186 38258
rect 66238 38206 66244 38258
rect 1576 37870 1582 37922
rect 1634 37870 1640 37922
rect 66180 37870 66186 37922
rect 66238 37870 66244 37922
rect 1576 37534 1582 37586
rect 1634 37534 1640 37586
rect 66180 37534 66186 37586
rect 66238 37534 66244 37586
rect 1576 37198 1582 37250
rect 1634 37198 1640 37250
rect 66180 37198 66186 37250
rect 66238 37198 66244 37250
rect 1576 36862 1582 36914
rect 1634 36862 1640 36914
rect 66180 36862 66186 36914
rect 66238 36862 66244 36914
rect 1576 36526 1582 36578
rect 1634 36526 1640 36578
rect 66180 36526 66186 36578
rect 66238 36526 66244 36578
rect 1576 36190 1582 36242
rect 1634 36190 1640 36242
rect 66180 36190 66186 36242
rect 66238 36190 66244 36242
rect 1576 35854 1582 35906
rect 1634 35854 1640 35906
rect 66180 35854 66186 35906
rect 66238 35854 66244 35906
rect 1576 35518 1582 35570
rect 1634 35518 1640 35570
rect 66180 35518 66186 35570
rect 66238 35518 66244 35570
rect 1576 35182 1582 35234
rect 1634 35182 1640 35234
rect 66180 35182 66186 35234
rect 66238 35182 66244 35234
rect 1576 34846 1582 34898
rect 1634 34846 1640 34898
rect 66180 34846 66186 34898
rect 66238 34846 66244 34898
rect 1576 34510 1582 34562
rect 1634 34510 1640 34562
rect 66180 34510 66186 34562
rect 66238 34510 66244 34562
rect 1576 34174 1582 34226
rect 1634 34174 1640 34226
rect 66180 34174 66186 34226
rect 66238 34174 66244 34226
rect 1576 33838 1582 33890
rect 1634 33838 1640 33890
rect 66180 33838 66186 33890
rect 66238 33838 66244 33890
rect 1576 33502 1582 33554
rect 1634 33502 1640 33554
rect 66180 33502 66186 33554
rect 66238 33502 66244 33554
rect 1576 33166 1582 33218
rect 1634 33166 1640 33218
rect 66180 33166 66186 33218
rect 66238 33166 66244 33218
rect 1576 32830 1582 32882
rect 1634 32830 1640 32882
rect 66180 32830 66186 32882
rect 66238 32830 66244 32882
rect 1576 32494 1582 32546
rect 1634 32494 1640 32546
rect 66180 32494 66186 32546
rect 66238 32494 66244 32546
rect 1576 32158 1582 32210
rect 1634 32158 1640 32210
rect 66180 32158 66186 32210
rect 66238 32158 66244 32210
rect 1576 31822 1582 31874
rect 1634 31822 1640 31874
rect 66180 31822 66186 31874
rect 66238 31822 66244 31874
rect 1576 31486 1582 31538
rect 1634 31486 1640 31538
rect 66180 31486 66186 31538
rect 66238 31486 66244 31538
rect 1576 31150 1582 31202
rect 1634 31150 1640 31202
rect 66180 31150 66186 31202
rect 66238 31150 66244 31202
rect 1576 30814 1582 30866
rect 1634 30814 1640 30866
rect 66180 30814 66186 30866
rect 66238 30814 66244 30866
rect 1576 30478 1582 30530
rect 1634 30478 1640 30530
rect 66180 30478 66186 30530
rect 66238 30478 66244 30530
rect 1576 30142 1582 30194
rect 1634 30142 1640 30194
rect 11405 30151 11411 30203
rect 11463 30151 11469 30203
rect 1576 29806 1582 29858
rect 1634 29806 1640 29858
rect 1576 29470 1582 29522
rect 1634 29470 1640 29522
rect 1576 29134 1582 29186
rect 1634 29134 1640 29186
rect 1576 28798 1582 28850
rect 1634 28798 1640 28850
rect 11325 28593 11331 28645
rect 11383 28593 11389 28645
rect 1576 28462 1582 28514
rect 1634 28462 1640 28514
rect 1576 28126 1582 28178
rect 1634 28126 1640 28178
rect 1576 27790 1582 27842
rect 1634 27790 1640 27842
rect 1576 27454 1582 27506
rect 1634 27454 1640 27506
rect 11245 27323 11251 27375
rect 11303 27323 11309 27375
rect 1576 27118 1582 27170
rect 1634 27118 1640 27170
rect 1576 26782 1582 26834
rect 1634 26782 1640 26834
rect 1576 26446 1582 26498
rect 1634 26446 1640 26498
rect 1576 26110 1582 26162
rect 1634 26110 1640 26162
rect 1576 25774 1582 25826
rect 1634 25774 1640 25826
rect 11165 25765 11171 25817
rect 11223 25765 11229 25817
rect 1576 25438 1582 25490
rect 1634 25438 1640 25490
rect 1576 25102 1582 25154
rect 1634 25102 1640 25154
rect 1576 24766 1582 24818
rect 1634 24766 1640 24818
rect 11085 24495 11091 24547
rect 11143 24495 11149 24547
rect 1576 24430 1582 24482
rect 1634 24430 1640 24482
rect 1576 24094 1582 24146
rect 1634 24094 1640 24146
rect 1576 23758 1582 23810
rect 1634 23758 1640 23810
rect 1576 23422 1582 23474
rect 1634 23422 1640 23474
rect 1576 23086 1582 23138
rect 1634 23086 1640 23138
rect 11005 22937 11011 22989
rect 11063 22937 11069 22989
rect 1576 22750 1582 22802
rect 1634 22750 1640 22802
rect 1576 22414 1582 22466
rect 1634 22414 1640 22466
rect 1576 22078 1582 22130
rect 1634 22078 1640 22130
rect 1576 21742 1582 21794
rect 1634 21742 1640 21794
rect 1576 21406 1582 21458
rect 1634 21406 1640 21458
rect 1576 21070 1582 21122
rect 1634 21070 1640 21122
rect 1576 20734 1582 20786
rect 1634 20734 1640 20786
rect 1576 20398 1582 20450
rect 1634 20398 1640 20450
rect 1576 20062 1582 20114
rect 1634 20062 1640 20114
rect 1576 19726 1582 19778
rect 1634 19726 1640 19778
rect 1576 19390 1582 19442
rect 1634 19390 1640 19442
rect 1576 19054 1582 19106
rect 1634 19054 1640 19106
rect 1576 18718 1582 18770
rect 1634 18718 1640 18770
rect 1576 18382 1582 18434
rect 1634 18382 1640 18434
rect 1576 18046 1582 18098
rect 1634 18046 1640 18098
rect 11023 17808 11051 22937
rect 11103 17808 11131 24495
rect 11183 17808 11211 25765
rect 11263 17808 11291 27323
rect 11343 17808 11371 28593
rect 11423 17808 11451 30151
rect 66180 30142 66186 30194
rect 66238 30142 66244 30194
rect 66180 29806 66186 29858
rect 66238 29806 66244 29858
rect 66180 29470 66186 29522
rect 66238 29470 66244 29522
rect 66180 29134 66186 29186
rect 66238 29134 66244 29186
rect 66180 28798 66186 28850
rect 66238 28798 66244 28850
rect 66180 28462 66186 28514
rect 66238 28462 66244 28514
rect 66180 28126 66186 28178
rect 66238 28126 66244 28178
rect 66180 27790 66186 27842
rect 66238 27790 66244 27842
rect 66180 27454 66186 27506
rect 66238 27454 66244 27506
rect 66180 27118 66186 27170
rect 66238 27118 66244 27170
rect 66180 26782 66186 26834
rect 66238 26782 66244 26834
rect 66180 26446 66186 26498
rect 66238 26446 66244 26498
rect 66180 26110 66186 26162
rect 66238 26110 66244 26162
rect 66180 25774 66186 25826
rect 66238 25774 66244 25826
rect 66180 25438 66186 25490
rect 66238 25438 66244 25490
rect 66180 25102 66186 25154
rect 66238 25102 66244 25154
rect 66180 24766 66186 24818
rect 66238 24766 66244 24818
rect 66180 24430 66186 24482
rect 66238 24430 66244 24482
rect 66180 24094 66186 24146
rect 66238 24094 66244 24146
rect 66180 23758 66186 23810
rect 66238 23758 66244 23810
rect 66180 23422 66186 23474
rect 66238 23422 66244 23474
rect 66180 23086 66186 23138
rect 66238 23086 66244 23138
rect 66180 22750 66186 22802
rect 66238 22750 66244 22802
rect 66180 22414 66186 22466
rect 66238 22414 66244 22466
rect 66180 22078 66186 22130
rect 66238 22078 66244 22130
rect 66180 21742 66186 21794
rect 66238 21742 66244 21794
rect 66180 21406 66186 21458
rect 66238 21406 66244 21458
rect 66180 21070 66186 21122
rect 66238 21070 66244 21122
rect 66180 20734 66186 20786
rect 66238 20734 66244 20786
rect 66180 20398 66186 20450
rect 66238 20398 66244 20450
rect 66180 20062 66186 20114
rect 66238 20062 66244 20114
rect 66180 19726 66186 19778
rect 66238 19726 66244 19778
rect 66180 19390 66186 19442
rect 66238 19390 66244 19442
rect 66180 19054 66186 19106
rect 66238 19054 66244 19106
rect 66180 18718 66186 18770
rect 66238 18718 66244 18770
rect 66180 18382 66186 18434
rect 66238 18382 66244 18434
rect 66180 18046 66186 18098
rect 66238 18046 66244 18098
rect 1576 17710 1582 17762
rect 1634 17710 1640 17762
rect 1576 17374 1582 17426
rect 1634 17374 1640 17426
rect 1576 17038 1582 17090
rect 1634 17038 1640 17090
rect 1576 16702 1582 16754
rect 1634 16702 1640 16754
rect 1576 16366 1582 16418
rect 1634 16366 1640 16418
rect 1576 16030 1582 16082
rect 1634 16030 1640 16082
rect 1576 15694 1582 15746
rect 1634 15694 1640 15746
rect 1576 15358 1582 15410
rect 1634 15358 1640 15410
rect 1576 15022 1582 15074
rect 1634 15022 1640 15074
rect 1576 14686 1582 14738
rect 1634 14686 1640 14738
rect 19016 14437 19022 14489
rect 19074 14437 19080 14489
rect 20907 14424 20913 14476
rect 20965 14424 20971 14476
rect 1576 14350 1582 14402
rect 1634 14350 1640 14402
rect 1576 14014 1582 14066
rect 1634 14014 1640 14066
rect 1576 13678 1582 13730
rect 1634 13678 1640 13730
rect 1576 13342 1582 13394
rect 1634 13342 1640 13394
rect 1576 13006 1582 13058
rect 1634 13006 1640 13058
rect 1576 12670 1582 12722
rect 1634 12670 1640 12722
rect 1576 12334 1582 12386
rect 1634 12334 1640 12386
rect 1576 11998 1582 12050
rect 1634 11998 1640 12050
rect 1576 11662 1582 11714
rect 1634 11662 1640 11714
rect 1576 11326 1582 11378
rect 1634 11326 1640 11378
rect 1576 10990 1582 11042
rect 1634 10990 1640 11042
rect 1576 10654 1582 10706
rect 1634 10654 1640 10706
rect 1576 10318 1582 10370
rect 1634 10318 1640 10370
rect 1576 9982 1582 10034
rect 1634 9982 1640 10034
rect 1576 9646 1582 9698
rect 1634 9646 1640 9698
rect 1576 9310 1582 9362
rect 1634 9310 1640 9362
rect 1576 8974 1582 9026
rect 1634 8974 1640 9026
rect 1576 8638 1582 8690
rect 1634 8638 1640 8690
rect 1576 8302 1582 8354
rect 1634 8302 1640 8354
rect 1576 7966 1582 8018
rect 1634 7966 1640 8018
rect 1576 7630 1582 7682
rect 1634 7630 1640 7682
rect 1576 7294 1582 7346
rect 1634 7294 1640 7346
rect 1576 6958 1582 7010
rect 1634 6958 1640 7010
rect 56285 6825 56313 17808
rect 56365 8383 56393 17808
rect 56445 9653 56473 17808
rect 56525 11211 56553 17808
rect 56605 12481 56633 17808
rect 56685 14039 56713 17808
rect 66180 17710 66186 17762
rect 66238 17710 66244 17762
rect 66180 17374 66186 17426
rect 66238 17374 66244 17426
rect 66180 17038 66186 17090
rect 66238 17038 66244 17090
rect 66180 16702 66186 16754
rect 66238 16702 66244 16754
rect 66180 16366 66186 16418
rect 66238 16366 66244 16418
rect 66180 16030 66186 16082
rect 66238 16030 66244 16082
rect 66180 15694 66186 15746
rect 66238 15694 66244 15746
rect 66180 15358 66186 15410
rect 66238 15358 66244 15410
rect 66180 15022 66186 15074
rect 66238 15022 66244 15074
rect 66180 14686 66186 14738
rect 66238 14686 66244 14738
rect 66180 14350 66186 14402
rect 66238 14350 66244 14402
rect 56667 13987 56673 14039
rect 56725 13987 56731 14039
rect 66180 14014 66186 14066
rect 66238 14014 66244 14066
rect 66180 13678 66186 13730
rect 66238 13678 66244 13730
rect 66180 13342 66186 13394
rect 66238 13342 66244 13394
rect 66180 13006 66186 13058
rect 66238 13006 66244 13058
rect 66180 12670 66186 12722
rect 66238 12670 66244 12722
rect 56587 12429 56593 12481
rect 56645 12429 56651 12481
rect 66180 12334 66186 12386
rect 66238 12334 66244 12386
rect 66180 11998 66186 12050
rect 66238 11998 66244 12050
rect 66180 11662 66186 11714
rect 66238 11662 66244 11714
rect 66180 11326 66186 11378
rect 66238 11326 66244 11378
rect 56507 11159 56513 11211
rect 56565 11159 56571 11211
rect 66180 10990 66186 11042
rect 66238 10990 66244 11042
rect 66180 10654 66186 10706
rect 66238 10654 66244 10706
rect 66180 10318 66186 10370
rect 66238 10318 66244 10370
rect 66180 9982 66186 10034
rect 66238 9982 66244 10034
rect 56427 9601 56433 9653
rect 56485 9601 56491 9653
rect 66180 9646 66186 9698
rect 66238 9646 66244 9698
rect 66180 9310 66186 9362
rect 66238 9310 66244 9362
rect 66180 8974 66186 9026
rect 66238 8974 66244 9026
rect 66180 8638 66186 8690
rect 66238 8638 66244 8690
rect 56347 8331 56353 8383
rect 56405 8331 56411 8383
rect 66180 8302 66186 8354
rect 66238 8302 66244 8354
rect 66180 7966 66186 8018
rect 66238 7966 66244 8018
rect 66180 7630 66186 7682
rect 66238 7630 66244 7682
rect 66180 7294 66186 7346
rect 66238 7294 66244 7346
rect 66180 6958 66186 7010
rect 66238 6958 66244 7010
rect 56267 6773 56273 6825
rect 56325 6773 56331 6825
rect 1576 6622 1582 6674
rect 1634 6622 1640 6674
rect 66180 6622 66186 6674
rect 66238 6622 66244 6674
rect 1576 6286 1582 6338
rect 1634 6286 1640 6338
rect 66180 6286 66186 6338
rect 66238 6286 66244 6338
rect 1576 5950 1582 6002
rect 1634 5950 1640 6002
rect 66180 5950 66186 6002
rect 66238 5950 66244 6002
rect 1576 5614 1582 5666
rect 1634 5614 1640 5666
rect 66180 5614 66186 5666
rect 66238 5614 66244 5666
rect 1576 5278 1582 5330
rect 1634 5278 1640 5330
rect 66180 5278 66186 5330
rect 66238 5278 66244 5330
rect 1576 4942 1582 4994
rect 1634 4942 1640 4994
rect 66180 4942 66186 4994
rect 66238 4942 66244 4994
rect 1576 4606 1582 4658
rect 1634 4606 1640 4658
rect 66180 4606 66186 4658
rect 66238 4606 66244 4658
rect 1576 4270 1582 4322
rect 1634 4270 1640 4322
rect 66180 4270 66186 4322
rect 66238 4270 66244 4322
rect 1576 3934 1582 3986
rect 1634 3934 1640 3986
rect 66180 3934 66186 3986
rect 66238 3934 66244 3986
rect 1576 3598 1582 3650
rect 1634 3598 1640 3650
rect 66180 3598 66186 3650
rect 66238 3598 66244 3650
rect 1576 3262 1582 3314
rect 1634 3262 1640 3314
rect 66180 3262 66186 3314
rect 66238 3262 66244 3314
rect 1576 2926 1582 2978
rect 1634 2926 1640 2978
rect 66180 2926 66186 2978
rect 66238 2926 66244 2978
rect 1576 2590 1582 2642
rect 1634 2590 1640 2642
rect 66180 2590 66186 2642
rect 66238 2590 66244 2642
rect 1576 2254 1582 2306
rect 1634 2254 1640 2306
rect 66180 2254 66186 2306
rect 66238 2254 66244 2306
rect 1576 1918 1582 1970
rect 1634 1918 1640 1970
rect 66180 1918 66186 1970
rect 66238 1918 66244 1970
rect 1496 1634 66324 1720
rect 1496 1582 1918 1634
rect 1970 1625 3598 1634
rect 3650 1625 5278 1634
rect 5330 1625 6958 1634
rect 7010 1625 8638 1634
rect 8690 1625 10318 1634
rect 10370 1625 11998 1634
rect 12050 1625 13678 1634
rect 13730 1625 15358 1634
rect 15410 1625 17038 1634
rect 17090 1625 18718 1634
rect 18770 1625 20398 1634
rect 20450 1625 22078 1634
rect 22130 1625 23758 1634
rect 23810 1625 25438 1634
rect 25490 1625 27118 1634
rect 27170 1625 28798 1634
rect 28850 1625 30478 1634
rect 30530 1625 32158 1634
rect 32210 1625 33838 1634
rect 33890 1625 35518 1634
rect 35570 1625 37198 1634
rect 37250 1625 38878 1634
rect 38930 1625 40558 1634
rect 40610 1625 42238 1634
rect 42290 1625 43918 1634
rect 43970 1625 45598 1634
rect 45650 1625 47278 1634
rect 47330 1625 48958 1634
rect 49010 1625 50638 1634
rect 50690 1625 52318 1634
rect 52370 1625 53998 1634
rect 54050 1625 55678 1634
rect 55730 1625 57358 1634
rect 57410 1625 59038 1634
rect 59090 1625 60718 1634
rect 60770 1625 62398 1634
rect 62450 1625 64078 1634
rect 64130 1625 65758 1634
rect 1970 1591 2263 1625
rect 2297 1591 2599 1625
rect 2633 1591 2935 1625
rect 2969 1591 3271 1625
rect 3305 1591 3598 1625
rect 3650 1591 3943 1625
rect 3977 1591 4279 1625
rect 4313 1591 4615 1625
rect 4649 1591 4951 1625
rect 4985 1591 5278 1625
rect 5330 1591 5623 1625
rect 5657 1591 5959 1625
rect 5993 1591 6295 1625
rect 6329 1591 6631 1625
rect 6665 1591 6958 1625
rect 7010 1591 7303 1625
rect 7337 1591 7639 1625
rect 7673 1591 7975 1625
rect 8009 1591 8311 1625
rect 8345 1591 8638 1625
rect 8690 1591 8983 1625
rect 9017 1591 9319 1625
rect 9353 1591 9655 1625
rect 9689 1591 9991 1625
rect 10025 1591 10318 1625
rect 10370 1591 10663 1625
rect 10697 1591 10999 1625
rect 11033 1591 11335 1625
rect 11369 1591 11671 1625
rect 11705 1591 11998 1625
rect 12050 1591 12343 1625
rect 12377 1591 12679 1625
rect 12713 1591 13015 1625
rect 13049 1591 13351 1625
rect 13385 1591 13678 1625
rect 13730 1591 14023 1625
rect 14057 1591 14359 1625
rect 14393 1591 14695 1625
rect 14729 1591 15031 1625
rect 15065 1591 15358 1625
rect 15410 1591 15703 1625
rect 15737 1591 16039 1625
rect 16073 1591 16375 1625
rect 16409 1591 16711 1625
rect 16745 1591 17038 1625
rect 17090 1591 17383 1625
rect 17417 1591 17719 1625
rect 17753 1591 18055 1625
rect 18089 1591 18391 1625
rect 18425 1591 18718 1625
rect 18770 1591 19063 1625
rect 19097 1591 19399 1625
rect 19433 1591 19735 1625
rect 19769 1591 20071 1625
rect 20105 1591 20398 1625
rect 20450 1591 20743 1625
rect 20777 1591 21079 1625
rect 21113 1591 21415 1625
rect 21449 1591 21751 1625
rect 21785 1591 22078 1625
rect 22130 1591 22423 1625
rect 22457 1591 22759 1625
rect 22793 1591 23095 1625
rect 23129 1591 23431 1625
rect 23465 1591 23758 1625
rect 23810 1591 24103 1625
rect 24137 1591 24439 1625
rect 24473 1591 24775 1625
rect 24809 1591 25111 1625
rect 25145 1591 25438 1625
rect 25490 1591 25783 1625
rect 25817 1591 26119 1625
rect 26153 1591 26455 1625
rect 26489 1591 26791 1625
rect 26825 1591 27118 1625
rect 27170 1591 27463 1625
rect 27497 1591 27799 1625
rect 27833 1591 28135 1625
rect 28169 1591 28471 1625
rect 28505 1591 28798 1625
rect 28850 1591 29143 1625
rect 29177 1591 29479 1625
rect 29513 1591 29815 1625
rect 29849 1591 30151 1625
rect 30185 1591 30478 1625
rect 30530 1591 30823 1625
rect 30857 1591 31159 1625
rect 31193 1591 31495 1625
rect 31529 1591 31831 1625
rect 31865 1591 32158 1625
rect 32210 1591 32503 1625
rect 32537 1591 32839 1625
rect 32873 1591 33175 1625
rect 33209 1591 33511 1625
rect 33545 1591 33838 1625
rect 33890 1591 34183 1625
rect 34217 1591 34519 1625
rect 34553 1591 34855 1625
rect 34889 1591 35191 1625
rect 35225 1591 35518 1625
rect 35570 1591 35863 1625
rect 35897 1591 36199 1625
rect 36233 1591 36535 1625
rect 36569 1591 36871 1625
rect 36905 1591 37198 1625
rect 37250 1591 37543 1625
rect 37577 1591 37879 1625
rect 37913 1591 38215 1625
rect 38249 1591 38551 1625
rect 38585 1591 38878 1625
rect 38930 1591 39223 1625
rect 39257 1591 39559 1625
rect 39593 1591 39895 1625
rect 39929 1591 40231 1625
rect 40265 1591 40558 1625
rect 40610 1591 40903 1625
rect 40937 1591 41239 1625
rect 41273 1591 41575 1625
rect 41609 1591 41911 1625
rect 41945 1591 42238 1625
rect 42290 1591 42583 1625
rect 42617 1591 42919 1625
rect 42953 1591 43255 1625
rect 43289 1591 43591 1625
rect 43625 1591 43918 1625
rect 43970 1591 44263 1625
rect 44297 1591 44599 1625
rect 44633 1591 44935 1625
rect 44969 1591 45271 1625
rect 45305 1591 45598 1625
rect 45650 1591 45943 1625
rect 45977 1591 46279 1625
rect 46313 1591 46615 1625
rect 46649 1591 46951 1625
rect 46985 1591 47278 1625
rect 47330 1591 47623 1625
rect 47657 1591 47959 1625
rect 47993 1591 48295 1625
rect 48329 1591 48631 1625
rect 48665 1591 48958 1625
rect 49010 1591 49303 1625
rect 49337 1591 49639 1625
rect 49673 1591 49975 1625
rect 50009 1591 50311 1625
rect 50345 1591 50638 1625
rect 50690 1591 50983 1625
rect 51017 1591 51319 1625
rect 51353 1591 51655 1625
rect 51689 1591 51991 1625
rect 52025 1591 52318 1625
rect 52370 1591 52663 1625
rect 52697 1591 52999 1625
rect 53033 1591 53335 1625
rect 53369 1591 53671 1625
rect 53705 1591 53998 1625
rect 54050 1591 54343 1625
rect 54377 1591 54679 1625
rect 54713 1591 55015 1625
rect 55049 1591 55351 1625
rect 55385 1591 55678 1625
rect 55730 1591 56023 1625
rect 56057 1591 56359 1625
rect 56393 1591 56695 1625
rect 56729 1591 57031 1625
rect 57065 1591 57358 1625
rect 57410 1591 57703 1625
rect 57737 1591 58039 1625
rect 58073 1591 58375 1625
rect 58409 1591 58711 1625
rect 58745 1591 59038 1625
rect 59090 1591 59383 1625
rect 59417 1591 59719 1625
rect 59753 1591 60055 1625
rect 60089 1591 60391 1625
rect 60425 1591 60718 1625
rect 60770 1591 61063 1625
rect 61097 1591 61399 1625
rect 61433 1591 61735 1625
rect 61769 1591 62071 1625
rect 62105 1591 62398 1625
rect 62450 1591 62743 1625
rect 62777 1591 63079 1625
rect 63113 1591 63415 1625
rect 63449 1591 63751 1625
rect 63785 1591 64078 1625
rect 64130 1591 64423 1625
rect 64457 1591 64759 1625
rect 64793 1591 65095 1625
rect 65129 1591 65431 1625
rect 65465 1591 65758 1625
rect 1970 1582 3598 1591
rect 3650 1582 5278 1591
rect 5330 1582 6958 1591
rect 7010 1582 8638 1591
rect 8690 1582 10318 1591
rect 10370 1582 11998 1591
rect 12050 1582 13678 1591
rect 13730 1582 15358 1591
rect 15410 1582 17038 1591
rect 17090 1582 18718 1591
rect 18770 1582 20398 1591
rect 20450 1582 22078 1591
rect 22130 1582 23758 1591
rect 23810 1582 25438 1591
rect 25490 1582 27118 1591
rect 27170 1582 28798 1591
rect 28850 1582 30478 1591
rect 30530 1582 32158 1591
rect 32210 1582 33838 1591
rect 33890 1582 35518 1591
rect 35570 1582 37198 1591
rect 37250 1582 38878 1591
rect 38930 1582 40558 1591
rect 40610 1582 42238 1591
rect 42290 1582 43918 1591
rect 43970 1582 45598 1591
rect 45650 1582 47278 1591
rect 47330 1582 48958 1591
rect 49010 1582 50638 1591
rect 50690 1582 52318 1591
rect 52370 1582 53998 1591
rect 54050 1582 55678 1591
rect 55730 1582 57358 1591
rect 57410 1582 59038 1591
rect 59090 1582 60718 1591
rect 60770 1582 62398 1591
rect 62450 1582 64078 1591
rect 64130 1582 65758 1591
rect 65810 1582 66324 1634
rect 1496 1496 66324 1582
<< via1 >>
rect 1918 51147 1970 51156
rect 3598 51147 3650 51156
rect 5278 51147 5330 51156
rect 6958 51147 7010 51156
rect 8638 51147 8690 51156
rect 10318 51147 10370 51156
rect 11998 51147 12050 51156
rect 13678 51147 13730 51156
rect 15358 51147 15410 51156
rect 17038 51147 17090 51156
rect 18718 51147 18770 51156
rect 20398 51147 20450 51156
rect 22078 51147 22130 51156
rect 23758 51147 23810 51156
rect 25438 51147 25490 51156
rect 27118 51147 27170 51156
rect 28798 51147 28850 51156
rect 30478 51147 30530 51156
rect 32158 51147 32210 51156
rect 33838 51147 33890 51156
rect 35518 51147 35570 51156
rect 37198 51147 37250 51156
rect 38878 51147 38930 51156
rect 40558 51147 40610 51156
rect 42238 51147 42290 51156
rect 43918 51147 43970 51156
rect 45598 51147 45650 51156
rect 47278 51147 47330 51156
rect 48958 51147 49010 51156
rect 50638 51147 50690 51156
rect 52318 51147 52370 51156
rect 53998 51147 54050 51156
rect 55678 51147 55730 51156
rect 57358 51147 57410 51156
rect 59038 51147 59090 51156
rect 60718 51147 60770 51156
rect 62398 51147 62450 51156
rect 64078 51147 64130 51156
rect 65758 51147 65810 51156
rect 1918 51113 1927 51147
rect 1927 51113 1961 51147
rect 1961 51113 1970 51147
rect 3598 51113 3607 51147
rect 3607 51113 3641 51147
rect 3641 51113 3650 51147
rect 5278 51113 5287 51147
rect 5287 51113 5321 51147
rect 5321 51113 5330 51147
rect 6958 51113 6967 51147
rect 6967 51113 7001 51147
rect 7001 51113 7010 51147
rect 8638 51113 8647 51147
rect 8647 51113 8681 51147
rect 8681 51113 8690 51147
rect 10318 51113 10327 51147
rect 10327 51113 10361 51147
rect 10361 51113 10370 51147
rect 11998 51113 12007 51147
rect 12007 51113 12041 51147
rect 12041 51113 12050 51147
rect 13678 51113 13687 51147
rect 13687 51113 13721 51147
rect 13721 51113 13730 51147
rect 15358 51113 15367 51147
rect 15367 51113 15401 51147
rect 15401 51113 15410 51147
rect 17038 51113 17047 51147
rect 17047 51113 17081 51147
rect 17081 51113 17090 51147
rect 18718 51113 18727 51147
rect 18727 51113 18761 51147
rect 18761 51113 18770 51147
rect 20398 51113 20407 51147
rect 20407 51113 20441 51147
rect 20441 51113 20450 51147
rect 22078 51113 22087 51147
rect 22087 51113 22121 51147
rect 22121 51113 22130 51147
rect 23758 51113 23767 51147
rect 23767 51113 23801 51147
rect 23801 51113 23810 51147
rect 25438 51113 25447 51147
rect 25447 51113 25481 51147
rect 25481 51113 25490 51147
rect 27118 51113 27127 51147
rect 27127 51113 27161 51147
rect 27161 51113 27170 51147
rect 28798 51113 28807 51147
rect 28807 51113 28841 51147
rect 28841 51113 28850 51147
rect 30478 51113 30487 51147
rect 30487 51113 30521 51147
rect 30521 51113 30530 51147
rect 32158 51113 32167 51147
rect 32167 51113 32201 51147
rect 32201 51113 32210 51147
rect 33838 51113 33847 51147
rect 33847 51113 33881 51147
rect 33881 51113 33890 51147
rect 35518 51113 35527 51147
rect 35527 51113 35561 51147
rect 35561 51113 35570 51147
rect 37198 51113 37207 51147
rect 37207 51113 37241 51147
rect 37241 51113 37250 51147
rect 38878 51113 38887 51147
rect 38887 51113 38921 51147
rect 38921 51113 38930 51147
rect 40558 51113 40567 51147
rect 40567 51113 40601 51147
rect 40601 51113 40610 51147
rect 42238 51113 42247 51147
rect 42247 51113 42281 51147
rect 42281 51113 42290 51147
rect 43918 51113 43927 51147
rect 43927 51113 43961 51147
rect 43961 51113 43970 51147
rect 45598 51113 45607 51147
rect 45607 51113 45641 51147
rect 45641 51113 45650 51147
rect 47278 51113 47287 51147
rect 47287 51113 47321 51147
rect 47321 51113 47330 51147
rect 48958 51113 48967 51147
rect 48967 51113 49001 51147
rect 49001 51113 49010 51147
rect 50638 51113 50647 51147
rect 50647 51113 50681 51147
rect 50681 51113 50690 51147
rect 52318 51113 52327 51147
rect 52327 51113 52361 51147
rect 52361 51113 52370 51147
rect 53998 51113 54007 51147
rect 54007 51113 54041 51147
rect 54041 51113 54050 51147
rect 55678 51113 55687 51147
rect 55687 51113 55721 51147
rect 55721 51113 55730 51147
rect 57358 51113 57367 51147
rect 57367 51113 57401 51147
rect 57401 51113 57410 51147
rect 59038 51113 59047 51147
rect 59047 51113 59081 51147
rect 59081 51113 59090 51147
rect 60718 51113 60727 51147
rect 60727 51113 60761 51147
rect 60761 51113 60770 51147
rect 62398 51113 62407 51147
rect 62407 51113 62441 51147
rect 62441 51113 62450 51147
rect 64078 51113 64087 51147
rect 64087 51113 64121 51147
rect 64121 51113 64130 51147
rect 65758 51113 65767 51147
rect 65767 51113 65801 51147
rect 65801 51113 65810 51147
rect 1918 51104 1970 51113
rect 3598 51104 3650 51113
rect 5278 51104 5330 51113
rect 6958 51104 7010 51113
rect 8638 51104 8690 51113
rect 10318 51104 10370 51113
rect 11998 51104 12050 51113
rect 13678 51104 13730 51113
rect 15358 51104 15410 51113
rect 17038 51104 17090 51113
rect 18718 51104 18770 51113
rect 20398 51104 20450 51113
rect 22078 51104 22130 51113
rect 23758 51104 23810 51113
rect 25438 51104 25490 51113
rect 27118 51104 27170 51113
rect 28798 51104 28850 51113
rect 30478 51104 30530 51113
rect 32158 51104 32210 51113
rect 33838 51104 33890 51113
rect 35518 51104 35570 51113
rect 37198 51104 37250 51113
rect 38878 51104 38930 51113
rect 40558 51104 40610 51113
rect 42238 51104 42290 51113
rect 43918 51104 43970 51113
rect 45598 51104 45650 51113
rect 47278 51104 47330 51113
rect 48958 51104 49010 51113
rect 50638 51104 50690 51113
rect 52318 51104 52370 51113
rect 53998 51104 54050 51113
rect 55678 51104 55730 51113
rect 57358 51104 57410 51113
rect 59038 51104 59090 51113
rect 60718 51104 60770 51113
rect 62398 51104 62450 51113
rect 64078 51104 64130 51113
rect 65758 51104 65810 51113
rect 1582 50681 1634 50690
rect 1582 50647 1591 50681
rect 1591 50647 1625 50681
rect 1625 50647 1634 50681
rect 1582 50638 1634 50647
rect 66186 50681 66238 50690
rect 66186 50647 66195 50681
rect 66195 50647 66229 50681
rect 66229 50647 66238 50681
rect 66186 50638 66238 50647
rect 1582 50345 1634 50354
rect 1582 50311 1591 50345
rect 1591 50311 1625 50345
rect 1625 50311 1634 50345
rect 1582 50302 1634 50311
rect 66186 50345 66238 50354
rect 66186 50311 66195 50345
rect 66195 50311 66229 50345
rect 66229 50311 66238 50345
rect 66186 50302 66238 50311
rect 1582 50009 1634 50018
rect 1582 49975 1591 50009
rect 1591 49975 1625 50009
rect 1625 49975 1634 50009
rect 1582 49966 1634 49975
rect 66186 50009 66238 50018
rect 66186 49975 66195 50009
rect 66195 49975 66229 50009
rect 66229 49975 66238 50009
rect 66186 49966 66238 49975
rect 1582 49673 1634 49682
rect 1582 49639 1591 49673
rect 1591 49639 1625 49673
rect 1625 49639 1634 49673
rect 1582 49630 1634 49639
rect 66186 49673 66238 49682
rect 66186 49639 66195 49673
rect 66195 49639 66229 49673
rect 66229 49639 66238 49673
rect 66186 49630 66238 49639
rect 1582 49337 1634 49346
rect 1582 49303 1591 49337
rect 1591 49303 1625 49337
rect 1625 49303 1634 49337
rect 1582 49294 1634 49303
rect 66186 49337 66238 49346
rect 66186 49303 66195 49337
rect 66195 49303 66229 49337
rect 66229 49303 66238 49337
rect 66186 49294 66238 49303
rect 1582 49001 1634 49010
rect 1582 48967 1591 49001
rect 1591 48967 1625 49001
rect 1625 48967 1634 49001
rect 1582 48958 1634 48967
rect 66186 49001 66238 49010
rect 66186 48967 66195 49001
rect 66195 48967 66229 49001
rect 66229 48967 66238 49001
rect 66186 48958 66238 48967
rect 1582 48665 1634 48674
rect 1582 48631 1591 48665
rect 1591 48631 1625 48665
rect 1625 48631 1634 48665
rect 1582 48622 1634 48631
rect 66186 48665 66238 48674
rect 66186 48631 66195 48665
rect 66195 48631 66229 48665
rect 66229 48631 66238 48665
rect 66186 48622 66238 48631
rect 1582 48329 1634 48338
rect 1582 48295 1591 48329
rect 1591 48295 1625 48329
rect 1625 48295 1634 48329
rect 1582 48286 1634 48295
rect 66186 48329 66238 48338
rect 66186 48295 66195 48329
rect 66195 48295 66229 48329
rect 66229 48295 66238 48329
rect 66186 48286 66238 48295
rect 1582 47993 1634 48002
rect 1582 47959 1591 47993
rect 1591 47959 1625 47993
rect 1625 47959 1634 47993
rect 1582 47950 1634 47959
rect 66186 47993 66238 48002
rect 66186 47959 66195 47993
rect 66195 47959 66229 47993
rect 66229 47959 66238 47993
rect 66186 47950 66238 47959
rect 1582 47657 1634 47666
rect 1582 47623 1591 47657
rect 1591 47623 1625 47657
rect 1625 47623 1634 47657
rect 1582 47614 1634 47623
rect 66186 47657 66238 47666
rect 66186 47623 66195 47657
rect 66195 47623 66229 47657
rect 66229 47623 66238 47657
rect 66186 47614 66238 47623
rect 1582 47321 1634 47330
rect 1582 47287 1591 47321
rect 1591 47287 1625 47321
rect 1625 47287 1634 47321
rect 1582 47278 1634 47287
rect 66186 47321 66238 47330
rect 66186 47287 66195 47321
rect 66195 47287 66229 47321
rect 66229 47287 66238 47321
rect 66186 47278 66238 47287
rect 1582 46985 1634 46994
rect 1582 46951 1591 46985
rect 1591 46951 1625 46985
rect 1625 46951 1634 46985
rect 1582 46942 1634 46951
rect 66186 46985 66238 46994
rect 66186 46951 66195 46985
rect 66195 46951 66229 46985
rect 66229 46951 66238 46985
rect 66186 46942 66238 46951
rect 23985 46835 24037 46887
rect 26481 46835 26533 46887
rect 28977 46835 29029 46887
rect 31473 46835 31525 46887
rect 33969 46835 34021 46887
rect 36465 46835 36517 46887
rect 38961 46835 39013 46887
rect 41457 46835 41509 46887
rect 1582 46649 1634 46658
rect 1582 46615 1591 46649
rect 1591 46615 1625 46649
rect 1625 46615 1634 46649
rect 1582 46606 1634 46615
rect 66186 46649 66238 46658
rect 66186 46615 66195 46649
rect 66195 46615 66229 46649
rect 66229 46615 66238 46649
rect 66186 46606 66238 46615
rect 1582 46313 1634 46322
rect 1582 46279 1591 46313
rect 1591 46279 1625 46313
rect 1625 46279 1634 46313
rect 1582 46270 1634 46279
rect 66186 46313 66238 46322
rect 66186 46279 66195 46313
rect 66195 46279 66229 46313
rect 66229 46279 66238 46313
rect 66186 46270 66238 46279
rect 1582 45977 1634 45986
rect 1582 45943 1591 45977
rect 1591 45943 1625 45977
rect 1625 45943 1634 45977
rect 1582 45934 1634 45943
rect 66186 45977 66238 45986
rect 66186 45943 66195 45977
rect 66195 45943 66229 45977
rect 66229 45943 66238 45977
rect 66186 45934 66238 45943
rect 1582 45641 1634 45650
rect 1582 45607 1591 45641
rect 1591 45607 1625 45641
rect 1625 45607 1634 45641
rect 1582 45598 1634 45607
rect 66186 45641 66238 45650
rect 66186 45607 66195 45641
rect 66195 45607 66229 45641
rect 66229 45607 66238 45641
rect 66186 45598 66238 45607
rect 1582 45305 1634 45314
rect 1582 45271 1591 45305
rect 1591 45271 1625 45305
rect 1625 45271 1634 45305
rect 1582 45262 1634 45271
rect 66186 45305 66238 45314
rect 66186 45271 66195 45305
rect 66195 45271 66229 45305
rect 66229 45271 66238 45305
rect 66186 45262 66238 45271
rect 1582 44969 1634 44978
rect 1582 44935 1591 44969
rect 1591 44935 1625 44969
rect 1625 44935 1634 44969
rect 1582 44926 1634 44935
rect 66186 44969 66238 44978
rect 66186 44935 66195 44969
rect 66195 44935 66229 44969
rect 66229 44935 66238 44969
rect 66186 44926 66238 44935
rect 1582 44633 1634 44642
rect 1582 44599 1591 44633
rect 1591 44599 1625 44633
rect 1625 44599 1634 44633
rect 1582 44590 1634 44599
rect 66186 44633 66238 44642
rect 66186 44599 66195 44633
rect 66195 44599 66229 44633
rect 66229 44599 66238 44633
rect 66186 44590 66238 44599
rect 1582 44297 1634 44306
rect 1582 44263 1591 44297
rect 1591 44263 1625 44297
rect 1625 44263 1634 44297
rect 1582 44254 1634 44263
rect 66186 44297 66238 44306
rect 66186 44263 66195 44297
rect 66195 44263 66229 44297
rect 66229 44263 66238 44297
rect 66186 44254 66238 44263
rect 1582 43961 1634 43970
rect 1582 43927 1591 43961
rect 1591 43927 1625 43961
rect 1625 43927 1634 43961
rect 1582 43918 1634 43927
rect 66186 43961 66238 43970
rect 66186 43927 66195 43961
rect 66195 43927 66229 43961
rect 66229 43927 66238 43961
rect 66186 43918 66238 43927
rect 1582 43625 1634 43634
rect 1582 43591 1591 43625
rect 1591 43591 1625 43625
rect 1625 43591 1634 43625
rect 1582 43582 1634 43591
rect 66186 43625 66238 43634
rect 66186 43591 66195 43625
rect 66195 43591 66229 43625
rect 66229 43591 66238 43625
rect 66186 43582 66238 43591
rect 1582 43289 1634 43298
rect 1582 43255 1591 43289
rect 1591 43255 1625 43289
rect 1625 43255 1634 43289
rect 1582 43246 1634 43255
rect 66186 43289 66238 43298
rect 66186 43255 66195 43289
rect 66195 43255 66229 43289
rect 66229 43255 66238 43289
rect 66186 43246 66238 43255
rect 1582 42953 1634 42962
rect 1582 42919 1591 42953
rect 1591 42919 1625 42953
rect 1625 42919 1634 42953
rect 1582 42910 1634 42919
rect 66186 42953 66238 42962
rect 66186 42919 66195 42953
rect 66195 42919 66229 42953
rect 66229 42919 66238 42953
rect 66186 42910 66238 42919
rect 1582 42617 1634 42626
rect 1582 42583 1591 42617
rect 1591 42583 1625 42617
rect 1625 42583 1634 42617
rect 1582 42574 1634 42583
rect 66186 42617 66238 42626
rect 66186 42583 66195 42617
rect 66195 42583 66229 42617
rect 66229 42583 66238 42617
rect 66186 42574 66238 42583
rect 1582 42281 1634 42290
rect 1582 42247 1591 42281
rect 1591 42247 1625 42281
rect 1625 42247 1634 42281
rect 1582 42238 1634 42247
rect 66186 42281 66238 42290
rect 66186 42247 66195 42281
rect 66195 42247 66229 42281
rect 66229 42247 66238 42281
rect 66186 42238 66238 42247
rect 1582 41945 1634 41954
rect 1582 41911 1591 41945
rect 1591 41911 1625 41945
rect 1625 41911 1634 41945
rect 1582 41902 1634 41911
rect 66186 41945 66238 41954
rect 66186 41911 66195 41945
rect 66195 41911 66229 41945
rect 66229 41911 66238 41945
rect 66186 41902 66238 41911
rect 1582 41609 1634 41618
rect 1582 41575 1591 41609
rect 1591 41575 1625 41609
rect 1625 41575 1634 41609
rect 1582 41566 1634 41575
rect 66186 41609 66238 41618
rect 66186 41575 66195 41609
rect 66195 41575 66229 41609
rect 66229 41575 66238 41609
rect 66186 41566 66238 41575
rect 1582 41273 1634 41282
rect 1582 41239 1591 41273
rect 1591 41239 1625 41273
rect 1625 41239 1634 41273
rect 1582 41230 1634 41239
rect 66186 41273 66238 41282
rect 66186 41239 66195 41273
rect 66195 41239 66229 41273
rect 66229 41239 66238 41273
rect 66186 41230 66238 41239
rect 1582 40937 1634 40946
rect 1582 40903 1591 40937
rect 1591 40903 1625 40937
rect 1625 40903 1634 40937
rect 1582 40894 1634 40903
rect 66186 40937 66238 40946
rect 66186 40903 66195 40937
rect 66195 40903 66229 40937
rect 66229 40903 66238 40937
rect 66186 40894 66238 40903
rect 1582 40601 1634 40610
rect 1582 40567 1591 40601
rect 1591 40567 1625 40601
rect 1625 40567 1634 40601
rect 1582 40558 1634 40567
rect 66186 40601 66238 40610
rect 66186 40567 66195 40601
rect 66195 40567 66229 40601
rect 66229 40567 66238 40601
rect 66186 40558 66238 40567
rect 1582 40265 1634 40274
rect 1582 40231 1591 40265
rect 1591 40231 1625 40265
rect 1625 40231 1634 40265
rect 1582 40222 1634 40231
rect 66186 40265 66238 40274
rect 66186 40231 66195 40265
rect 66195 40231 66229 40265
rect 66229 40231 66238 40265
rect 66186 40222 66238 40231
rect 46771 40100 46823 40152
rect 48662 40087 48714 40139
rect 1582 39929 1634 39938
rect 1582 39895 1591 39929
rect 1591 39895 1625 39929
rect 1625 39895 1634 39929
rect 1582 39886 1634 39895
rect 66186 39929 66238 39938
rect 66186 39895 66195 39929
rect 66195 39895 66229 39929
rect 66229 39895 66238 39929
rect 66186 39886 66238 39895
rect 1582 39593 1634 39602
rect 1582 39559 1591 39593
rect 1591 39559 1625 39593
rect 1625 39559 1634 39593
rect 1582 39550 1634 39559
rect 66186 39593 66238 39602
rect 66186 39559 66195 39593
rect 66195 39559 66229 39593
rect 66229 39559 66238 39593
rect 66186 39550 66238 39559
rect 1582 39257 1634 39266
rect 1582 39223 1591 39257
rect 1591 39223 1625 39257
rect 1625 39223 1634 39257
rect 1582 39214 1634 39223
rect 66186 39257 66238 39266
rect 66186 39223 66195 39257
rect 66195 39223 66229 39257
rect 66229 39223 66238 39257
rect 66186 39214 66238 39223
rect 1582 38921 1634 38930
rect 1582 38887 1591 38921
rect 1591 38887 1625 38921
rect 1625 38887 1634 38921
rect 1582 38878 1634 38887
rect 66186 38921 66238 38930
rect 66186 38887 66195 38921
rect 66195 38887 66229 38921
rect 66229 38887 66238 38921
rect 66186 38878 66238 38887
rect 1582 38585 1634 38594
rect 1582 38551 1591 38585
rect 1591 38551 1625 38585
rect 1625 38551 1634 38585
rect 1582 38542 1634 38551
rect 66186 38585 66238 38594
rect 66186 38551 66195 38585
rect 66195 38551 66229 38585
rect 66229 38551 66238 38585
rect 66186 38542 66238 38551
rect 1582 38249 1634 38258
rect 1582 38215 1591 38249
rect 1591 38215 1625 38249
rect 1625 38215 1634 38249
rect 1582 38206 1634 38215
rect 66186 38249 66238 38258
rect 66186 38215 66195 38249
rect 66195 38215 66229 38249
rect 66229 38215 66238 38249
rect 66186 38206 66238 38215
rect 1582 37913 1634 37922
rect 1582 37879 1591 37913
rect 1591 37879 1625 37913
rect 1625 37879 1634 37913
rect 1582 37870 1634 37879
rect 66186 37913 66238 37922
rect 66186 37879 66195 37913
rect 66195 37879 66229 37913
rect 66229 37879 66238 37913
rect 66186 37870 66238 37879
rect 1582 37577 1634 37586
rect 1582 37543 1591 37577
rect 1591 37543 1625 37577
rect 1625 37543 1634 37577
rect 1582 37534 1634 37543
rect 66186 37577 66238 37586
rect 66186 37543 66195 37577
rect 66195 37543 66229 37577
rect 66229 37543 66238 37577
rect 66186 37534 66238 37543
rect 1582 37241 1634 37250
rect 1582 37207 1591 37241
rect 1591 37207 1625 37241
rect 1625 37207 1634 37241
rect 1582 37198 1634 37207
rect 66186 37241 66238 37250
rect 66186 37207 66195 37241
rect 66195 37207 66229 37241
rect 66229 37207 66238 37241
rect 66186 37198 66238 37207
rect 1582 36905 1634 36914
rect 1582 36871 1591 36905
rect 1591 36871 1625 36905
rect 1625 36871 1634 36905
rect 1582 36862 1634 36871
rect 66186 36905 66238 36914
rect 66186 36871 66195 36905
rect 66195 36871 66229 36905
rect 66229 36871 66238 36905
rect 66186 36862 66238 36871
rect 1582 36569 1634 36578
rect 1582 36535 1591 36569
rect 1591 36535 1625 36569
rect 1625 36535 1634 36569
rect 1582 36526 1634 36535
rect 66186 36569 66238 36578
rect 66186 36535 66195 36569
rect 66195 36535 66229 36569
rect 66229 36535 66238 36569
rect 66186 36526 66238 36535
rect 1582 36233 1634 36242
rect 1582 36199 1591 36233
rect 1591 36199 1625 36233
rect 1625 36199 1634 36233
rect 1582 36190 1634 36199
rect 66186 36233 66238 36242
rect 66186 36199 66195 36233
rect 66195 36199 66229 36233
rect 66229 36199 66238 36233
rect 66186 36190 66238 36199
rect 1582 35897 1634 35906
rect 1582 35863 1591 35897
rect 1591 35863 1625 35897
rect 1625 35863 1634 35897
rect 1582 35854 1634 35863
rect 66186 35897 66238 35906
rect 66186 35863 66195 35897
rect 66195 35863 66229 35897
rect 66229 35863 66238 35897
rect 66186 35854 66238 35863
rect 1582 35561 1634 35570
rect 1582 35527 1591 35561
rect 1591 35527 1625 35561
rect 1625 35527 1634 35561
rect 1582 35518 1634 35527
rect 66186 35561 66238 35570
rect 66186 35527 66195 35561
rect 66195 35527 66229 35561
rect 66229 35527 66238 35561
rect 66186 35518 66238 35527
rect 1582 35225 1634 35234
rect 1582 35191 1591 35225
rect 1591 35191 1625 35225
rect 1625 35191 1634 35225
rect 1582 35182 1634 35191
rect 66186 35225 66238 35234
rect 66186 35191 66195 35225
rect 66195 35191 66229 35225
rect 66229 35191 66238 35225
rect 66186 35182 66238 35191
rect 1582 34889 1634 34898
rect 1582 34855 1591 34889
rect 1591 34855 1625 34889
rect 1625 34855 1634 34889
rect 1582 34846 1634 34855
rect 66186 34889 66238 34898
rect 66186 34855 66195 34889
rect 66195 34855 66229 34889
rect 66229 34855 66238 34889
rect 66186 34846 66238 34855
rect 1582 34553 1634 34562
rect 1582 34519 1591 34553
rect 1591 34519 1625 34553
rect 1625 34519 1634 34553
rect 1582 34510 1634 34519
rect 66186 34553 66238 34562
rect 66186 34519 66195 34553
rect 66195 34519 66229 34553
rect 66229 34519 66238 34553
rect 66186 34510 66238 34519
rect 1582 34217 1634 34226
rect 1582 34183 1591 34217
rect 1591 34183 1625 34217
rect 1625 34183 1634 34217
rect 1582 34174 1634 34183
rect 66186 34217 66238 34226
rect 66186 34183 66195 34217
rect 66195 34183 66229 34217
rect 66229 34183 66238 34217
rect 66186 34174 66238 34183
rect 1582 33881 1634 33890
rect 1582 33847 1591 33881
rect 1591 33847 1625 33881
rect 1625 33847 1634 33881
rect 1582 33838 1634 33847
rect 66186 33881 66238 33890
rect 66186 33847 66195 33881
rect 66195 33847 66229 33881
rect 66229 33847 66238 33881
rect 66186 33838 66238 33847
rect 1582 33545 1634 33554
rect 1582 33511 1591 33545
rect 1591 33511 1625 33545
rect 1625 33511 1634 33545
rect 1582 33502 1634 33511
rect 66186 33545 66238 33554
rect 66186 33511 66195 33545
rect 66195 33511 66229 33545
rect 66229 33511 66238 33545
rect 66186 33502 66238 33511
rect 1582 33209 1634 33218
rect 1582 33175 1591 33209
rect 1591 33175 1625 33209
rect 1625 33175 1634 33209
rect 1582 33166 1634 33175
rect 66186 33209 66238 33218
rect 66186 33175 66195 33209
rect 66195 33175 66229 33209
rect 66229 33175 66238 33209
rect 66186 33166 66238 33175
rect 1582 32873 1634 32882
rect 1582 32839 1591 32873
rect 1591 32839 1625 32873
rect 1625 32839 1634 32873
rect 1582 32830 1634 32839
rect 66186 32873 66238 32882
rect 66186 32839 66195 32873
rect 66195 32839 66229 32873
rect 66229 32839 66238 32873
rect 66186 32830 66238 32839
rect 1582 32537 1634 32546
rect 1582 32503 1591 32537
rect 1591 32503 1625 32537
rect 1625 32503 1634 32537
rect 1582 32494 1634 32503
rect 66186 32537 66238 32546
rect 66186 32503 66195 32537
rect 66195 32503 66229 32537
rect 66229 32503 66238 32537
rect 66186 32494 66238 32503
rect 1582 32201 1634 32210
rect 1582 32167 1591 32201
rect 1591 32167 1625 32201
rect 1625 32167 1634 32201
rect 1582 32158 1634 32167
rect 66186 32201 66238 32210
rect 66186 32167 66195 32201
rect 66195 32167 66229 32201
rect 66229 32167 66238 32201
rect 66186 32158 66238 32167
rect 1582 31865 1634 31874
rect 1582 31831 1591 31865
rect 1591 31831 1625 31865
rect 1625 31831 1634 31865
rect 1582 31822 1634 31831
rect 66186 31865 66238 31874
rect 66186 31831 66195 31865
rect 66195 31831 66229 31865
rect 66229 31831 66238 31865
rect 66186 31822 66238 31831
rect 1582 31529 1634 31538
rect 1582 31495 1591 31529
rect 1591 31495 1625 31529
rect 1625 31495 1634 31529
rect 1582 31486 1634 31495
rect 66186 31529 66238 31538
rect 66186 31495 66195 31529
rect 66195 31495 66229 31529
rect 66229 31495 66238 31529
rect 66186 31486 66238 31495
rect 1582 31193 1634 31202
rect 1582 31159 1591 31193
rect 1591 31159 1625 31193
rect 1625 31159 1634 31193
rect 1582 31150 1634 31159
rect 66186 31193 66238 31202
rect 66186 31159 66195 31193
rect 66195 31159 66229 31193
rect 66229 31159 66238 31193
rect 66186 31150 66238 31159
rect 1582 30857 1634 30866
rect 1582 30823 1591 30857
rect 1591 30823 1625 30857
rect 1625 30823 1634 30857
rect 1582 30814 1634 30823
rect 66186 30857 66238 30866
rect 66186 30823 66195 30857
rect 66195 30823 66229 30857
rect 66229 30823 66238 30857
rect 66186 30814 66238 30823
rect 1582 30521 1634 30530
rect 1582 30487 1591 30521
rect 1591 30487 1625 30521
rect 1625 30487 1634 30521
rect 1582 30478 1634 30487
rect 66186 30521 66238 30530
rect 66186 30487 66195 30521
rect 66195 30487 66229 30521
rect 66229 30487 66238 30521
rect 66186 30478 66238 30487
rect 1582 30185 1634 30194
rect 1582 30151 1591 30185
rect 1591 30151 1625 30185
rect 1625 30151 1634 30185
rect 1582 30142 1634 30151
rect 11411 30151 11463 30203
rect 1582 29849 1634 29858
rect 1582 29815 1591 29849
rect 1591 29815 1625 29849
rect 1625 29815 1634 29849
rect 1582 29806 1634 29815
rect 1582 29513 1634 29522
rect 1582 29479 1591 29513
rect 1591 29479 1625 29513
rect 1625 29479 1634 29513
rect 1582 29470 1634 29479
rect 1582 29177 1634 29186
rect 1582 29143 1591 29177
rect 1591 29143 1625 29177
rect 1625 29143 1634 29177
rect 1582 29134 1634 29143
rect 1582 28841 1634 28850
rect 1582 28807 1591 28841
rect 1591 28807 1625 28841
rect 1625 28807 1634 28841
rect 1582 28798 1634 28807
rect 11331 28593 11383 28645
rect 1582 28505 1634 28514
rect 1582 28471 1591 28505
rect 1591 28471 1625 28505
rect 1625 28471 1634 28505
rect 1582 28462 1634 28471
rect 1582 28169 1634 28178
rect 1582 28135 1591 28169
rect 1591 28135 1625 28169
rect 1625 28135 1634 28169
rect 1582 28126 1634 28135
rect 1582 27833 1634 27842
rect 1582 27799 1591 27833
rect 1591 27799 1625 27833
rect 1625 27799 1634 27833
rect 1582 27790 1634 27799
rect 1582 27497 1634 27506
rect 1582 27463 1591 27497
rect 1591 27463 1625 27497
rect 1625 27463 1634 27497
rect 1582 27454 1634 27463
rect 11251 27323 11303 27375
rect 1582 27161 1634 27170
rect 1582 27127 1591 27161
rect 1591 27127 1625 27161
rect 1625 27127 1634 27161
rect 1582 27118 1634 27127
rect 1582 26825 1634 26834
rect 1582 26791 1591 26825
rect 1591 26791 1625 26825
rect 1625 26791 1634 26825
rect 1582 26782 1634 26791
rect 1582 26489 1634 26498
rect 1582 26455 1591 26489
rect 1591 26455 1625 26489
rect 1625 26455 1634 26489
rect 1582 26446 1634 26455
rect 1582 26153 1634 26162
rect 1582 26119 1591 26153
rect 1591 26119 1625 26153
rect 1625 26119 1634 26153
rect 1582 26110 1634 26119
rect 1582 25817 1634 25826
rect 1582 25783 1591 25817
rect 1591 25783 1625 25817
rect 1625 25783 1634 25817
rect 1582 25774 1634 25783
rect 11171 25765 11223 25817
rect 1582 25481 1634 25490
rect 1582 25447 1591 25481
rect 1591 25447 1625 25481
rect 1625 25447 1634 25481
rect 1582 25438 1634 25447
rect 1582 25145 1634 25154
rect 1582 25111 1591 25145
rect 1591 25111 1625 25145
rect 1625 25111 1634 25145
rect 1582 25102 1634 25111
rect 1582 24809 1634 24818
rect 1582 24775 1591 24809
rect 1591 24775 1625 24809
rect 1625 24775 1634 24809
rect 1582 24766 1634 24775
rect 11091 24495 11143 24547
rect 1582 24473 1634 24482
rect 1582 24439 1591 24473
rect 1591 24439 1625 24473
rect 1625 24439 1634 24473
rect 1582 24430 1634 24439
rect 1582 24137 1634 24146
rect 1582 24103 1591 24137
rect 1591 24103 1625 24137
rect 1625 24103 1634 24137
rect 1582 24094 1634 24103
rect 1582 23801 1634 23810
rect 1582 23767 1591 23801
rect 1591 23767 1625 23801
rect 1625 23767 1634 23801
rect 1582 23758 1634 23767
rect 1582 23465 1634 23474
rect 1582 23431 1591 23465
rect 1591 23431 1625 23465
rect 1625 23431 1634 23465
rect 1582 23422 1634 23431
rect 1582 23129 1634 23138
rect 1582 23095 1591 23129
rect 1591 23095 1625 23129
rect 1625 23095 1634 23129
rect 1582 23086 1634 23095
rect 11011 22937 11063 22989
rect 1582 22793 1634 22802
rect 1582 22759 1591 22793
rect 1591 22759 1625 22793
rect 1625 22759 1634 22793
rect 1582 22750 1634 22759
rect 1582 22457 1634 22466
rect 1582 22423 1591 22457
rect 1591 22423 1625 22457
rect 1625 22423 1634 22457
rect 1582 22414 1634 22423
rect 1582 22121 1634 22130
rect 1582 22087 1591 22121
rect 1591 22087 1625 22121
rect 1625 22087 1634 22121
rect 1582 22078 1634 22087
rect 1582 21785 1634 21794
rect 1582 21751 1591 21785
rect 1591 21751 1625 21785
rect 1625 21751 1634 21785
rect 1582 21742 1634 21751
rect 1582 21449 1634 21458
rect 1582 21415 1591 21449
rect 1591 21415 1625 21449
rect 1625 21415 1634 21449
rect 1582 21406 1634 21415
rect 1582 21113 1634 21122
rect 1582 21079 1591 21113
rect 1591 21079 1625 21113
rect 1625 21079 1634 21113
rect 1582 21070 1634 21079
rect 1582 20777 1634 20786
rect 1582 20743 1591 20777
rect 1591 20743 1625 20777
rect 1625 20743 1634 20777
rect 1582 20734 1634 20743
rect 1582 20441 1634 20450
rect 1582 20407 1591 20441
rect 1591 20407 1625 20441
rect 1625 20407 1634 20441
rect 1582 20398 1634 20407
rect 1582 20105 1634 20114
rect 1582 20071 1591 20105
rect 1591 20071 1625 20105
rect 1625 20071 1634 20105
rect 1582 20062 1634 20071
rect 1582 19769 1634 19778
rect 1582 19735 1591 19769
rect 1591 19735 1625 19769
rect 1625 19735 1634 19769
rect 1582 19726 1634 19735
rect 1582 19433 1634 19442
rect 1582 19399 1591 19433
rect 1591 19399 1625 19433
rect 1625 19399 1634 19433
rect 1582 19390 1634 19399
rect 1582 19097 1634 19106
rect 1582 19063 1591 19097
rect 1591 19063 1625 19097
rect 1625 19063 1634 19097
rect 1582 19054 1634 19063
rect 1582 18761 1634 18770
rect 1582 18727 1591 18761
rect 1591 18727 1625 18761
rect 1625 18727 1634 18761
rect 1582 18718 1634 18727
rect 1582 18425 1634 18434
rect 1582 18391 1591 18425
rect 1591 18391 1625 18425
rect 1625 18391 1634 18425
rect 1582 18382 1634 18391
rect 1582 18089 1634 18098
rect 1582 18055 1591 18089
rect 1591 18055 1625 18089
rect 1625 18055 1634 18089
rect 1582 18046 1634 18055
rect 66186 30185 66238 30194
rect 66186 30151 66195 30185
rect 66195 30151 66229 30185
rect 66229 30151 66238 30185
rect 66186 30142 66238 30151
rect 66186 29849 66238 29858
rect 66186 29815 66195 29849
rect 66195 29815 66229 29849
rect 66229 29815 66238 29849
rect 66186 29806 66238 29815
rect 66186 29513 66238 29522
rect 66186 29479 66195 29513
rect 66195 29479 66229 29513
rect 66229 29479 66238 29513
rect 66186 29470 66238 29479
rect 66186 29177 66238 29186
rect 66186 29143 66195 29177
rect 66195 29143 66229 29177
rect 66229 29143 66238 29177
rect 66186 29134 66238 29143
rect 66186 28841 66238 28850
rect 66186 28807 66195 28841
rect 66195 28807 66229 28841
rect 66229 28807 66238 28841
rect 66186 28798 66238 28807
rect 66186 28505 66238 28514
rect 66186 28471 66195 28505
rect 66195 28471 66229 28505
rect 66229 28471 66238 28505
rect 66186 28462 66238 28471
rect 66186 28169 66238 28178
rect 66186 28135 66195 28169
rect 66195 28135 66229 28169
rect 66229 28135 66238 28169
rect 66186 28126 66238 28135
rect 66186 27833 66238 27842
rect 66186 27799 66195 27833
rect 66195 27799 66229 27833
rect 66229 27799 66238 27833
rect 66186 27790 66238 27799
rect 66186 27497 66238 27506
rect 66186 27463 66195 27497
rect 66195 27463 66229 27497
rect 66229 27463 66238 27497
rect 66186 27454 66238 27463
rect 66186 27161 66238 27170
rect 66186 27127 66195 27161
rect 66195 27127 66229 27161
rect 66229 27127 66238 27161
rect 66186 27118 66238 27127
rect 66186 26825 66238 26834
rect 66186 26791 66195 26825
rect 66195 26791 66229 26825
rect 66229 26791 66238 26825
rect 66186 26782 66238 26791
rect 66186 26489 66238 26498
rect 66186 26455 66195 26489
rect 66195 26455 66229 26489
rect 66229 26455 66238 26489
rect 66186 26446 66238 26455
rect 66186 26153 66238 26162
rect 66186 26119 66195 26153
rect 66195 26119 66229 26153
rect 66229 26119 66238 26153
rect 66186 26110 66238 26119
rect 66186 25817 66238 25826
rect 66186 25783 66195 25817
rect 66195 25783 66229 25817
rect 66229 25783 66238 25817
rect 66186 25774 66238 25783
rect 66186 25481 66238 25490
rect 66186 25447 66195 25481
rect 66195 25447 66229 25481
rect 66229 25447 66238 25481
rect 66186 25438 66238 25447
rect 66186 25145 66238 25154
rect 66186 25111 66195 25145
rect 66195 25111 66229 25145
rect 66229 25111 66238 25145
rect 66186 25102 66238 25111
rect 66186 24809 66238 24818
rect 66186 24775 66195 24809
rect 66195 24775 66229 24809
rect 66229 24775 66238 24809
rect 66186 24766 66238 24775
rect 66186 24473 66238 24482
rect 66186 24439 66195 24473
rect 66195 24439 66229 24473
rect 66229 24439 66238 24473
rect 66186 24430 66238 24439
rect 66186 24137 66238 24146
rect 66186 24103 66195 24137
rect 66195 24103 66229 24137
rect 66229 24103 66238 24137
rect 66186 24094 66238 24103
rect 66186 23801 66238 23810
rect 66186 23767 66195 23801
rect 66195 23767 66229 23801
rect 66229 23767 66238 23801
rect 66186 23758 66238 23767
rect 66186 23465 66238 23474
rect 66186 23431 66195 23465
rect 66195 23431 66229 23465
rect 66229 23431 66238 23465
rect 66186 23422 66238 23431
rect 66186 23129 66238 23138
rect 66186 23095 66195 23129
rect 66195 23095 66229 23129
rect 66229 23095 66238 23129
rect 66186 23086 66238 23095
rect 66186 22793 66238 22802
rect 66186 22759 66195 22793
rect 66195 22759 66229 22793
rect 66229 22759 66238 22793
rect 66186 22750 66238 22759
rect 66186 22457 66238 22466
rect 66186 22423 66195 22457
rect 66195 22423 66229 22457
rect 66229 22423 66238 22457
rect 66186 22414 66238 22423
rect 66186 22121 66238 22130
rect 66186 22087 66195 22121
rect 66195 22087 66229 22121
rect 66229 22087 66238 22121
rect 66186 22078 66238 22087
rect 66186 21785 66238 21794
rect 66186 21751 66195 21785
rect 66195 21751 66229 21785
rect 66229 21751 66238 21785
rect 66186 21742 66238 21751
rect 66186 21449 66238 21458
rect 66186 21415 66195 21449
rect 66195 21415 66229 21449
rect 66229 21415 66238 21449
rect 66186 21406 66238 21415
rect 66186 21113 66238 21122
rect 66186 21079 66195 21113
rect 66195 21079 66229 21113
rect 66229 21079 66238 21113
rect 66186 21070 66238 21079
rect 66186 20777 66238 20786
rect 66186 20743 66195 20777
rect 66195 20743 66229 20777
rect 66229 20743 66238 20777
rect 66186 20734 66238 20743
rect 66186 20441 66238 20450
rect 66186 20407 66195 20441
rect 66195 20407 66229 20441
rect 66229 20407 66238 20441
rect 66186 20398 66238 20407
rect 66186 20105 66238 20114
rect 66186 20071 66195 20105
rect 66195 20071 66229 20105
rect 66229 20071 66238 20105
rect 66186 20062 66238 20071
rect 66186 19769 66238 19778
rect 66186 19735 66195 19769
rect 66195 19735 66229 19769
rect 66229 19735 66238 19769
rect 66186 19726 66238 19735
rect 66186 19433 66238 19442
rect 66186 19399 66195 19433
rect 66195 19399 66229 19433
rect 66229 19399 66238 19433
rect 66186 19390 66238 19399
rect 66186 19097 66238 19106
rect 66186 19063 66195 19097
rect 66195 19063 66229 19097
rect 66229 19063 66238 19097
rect 66186 19054 66238 19063
rect 66186 18761 66238 18770
rect 66186 18727 66195 18761
rect 66195 18727 66229 18761
rect 66229 18727 66238 18761
rect 66186 18718 66238 18727
rect 66186 18425 66238 18434
rect 66186 18391 66195 18425
rect 66195 18391 66229 18425
rect 66229 18391 66238 18425
rect 66186 18382 66238 18391
rect 66186 18089 66238 18098
rect 66186 18055 66195 18089
rect 66195 18055 66229 18089
rect 66229 18055 66238 18089
rect 66186 18046 66238 18055
rect 1582 17753 1634 17762
rect 1582 17719 1591 17753
rect 1591 17719 1625 17753
rect 1625 17719 1634 17753
rect 1582 17710 1634 17719
rect 1582 17417 1634 17426
rect 1582 17383 1591 17417
rect 1591 17383 1625 17417
rect 1625 17383 1634 17417
rect 1582 17374 1634 17383
rect 1582 17081 1634 17090
rect 1582 17047 1591 17081
rect 1591 17047 1625 17081
rect 1625 17047 1634 17081
rect 1582 17038 1634 17047
rect 1582 16745 1634 16754
rect 1582 16711 1591 16745
rect 1591 16711 1625 16745
rect 1625 16711 1634 16745
rect 1582 16702 1634 16711
rect 1582 16409 1634 16418
rect 1582 16375 1591 16409
rect 1591 16375 1625 16409
rect 1625 16375 1634 16409
rect 1582 16366 1634 16375
rect 1582 16073 1634 16082
rect 1582 16039 1591 16073
rect 1591 16039 1625 16073
rect 1625 16039 1634 16073
rect 1582 16030 1634 16039
rect 1582 15737 1634 15746
rect 1582 15703 1591 15737
rect 1591 15703 1625 15737
rect 1625 15703 1634 15737
rect 1582 15694 1634 15703
rect 1582 15401 1634 15410
rect 1582 15367 1591 15401
rect 1591 15367 1625 15401
rect 1625 15367 1634 15401
rect 1582 15358 1634 15367
rect 1582 15065 1634 15074
rect 1582 15031 1591 15065
rect 1591 15031 1625 15065
rect 1625 15031 1634 15065
rect 1582 15022 1634 15031
rect 1582 14729 1634 14738
rect 1582 14695 1591 14729
rect 1591 14695 1625 14729
rect 1625 14695 1634 14729
rect 1582 14686 1634 14695
rect 19022 14437 19074 14489
rect 20913 14424 20965 14476
rect 1582 14393 1634 14402
rect 1582 14359 1591 14393
rect 1591 14359 1625 14393
rect 1625 14359 1634 14393
rect 1582 14350 1634 14359
rect 1582 14057 1634 14066
rect 1582 14023 1591 14057
rect 1591 14023 1625 14057
rect 1625 14023 1634 14057
rect 1582 14014 1634 14023
rect 1582 13721 1634 13730
rect 1582 13687 1591 13721
rect 1591 13687 1625 13721
rect 1625 13687 1634 13721
rect 1582 13678 1634 13687
rect 1582 13385 1634 13394
rect 1582 13351 1591 13385
rect 1591 13351 1625 13385
rect 1625 13351 1634 13385
rect 1582 13342 1634 13351
rect 1582 13049 1634 13058
rect 1582 13015 1591 13049
rect 1591 13015 1625 13049
rect 1625 13015 1634 13049
rect 1582 13006 1634 13015
rect 1582 12713 1634 12722
rect 1582 12679 1591 12713
rect 1591 12679 1625 12713
rect 1625 12679 1634 12713
rect 1582 12670 1634 12679
rect 1582 12377 1634 12386
rect 1582 12343 1591 12377
rect 1591 12343 1625 12377
rect 1625 12343 1634 12377
rect 1582 12334 1634 12343
rect 1582 12041 1634 12050
rect 1582 12007 1591 12041
rect 1591 12007 1625 12041
rect 1625 12007 1634 12041
rect 1582 11998 1634 12007
rect 1582 11705 1634 11714
rect 1582 11671 1591 11705
rect 1591 11671 1625 11705
rect 1625 11671 1634 11705
rect 1582 11662 1634 11671
rect 1582 11369 1634 11378
rect 1582 11335 1591 11369
rect 1591 11335 1625 11369
rect 1625 11335 1634 11369
rect 1582 11326 1634 11335
rect 1582 11033 1634 11042
rect 1582 10999 1591 11033
rect 1591 10999 1625 11033
rect 1625 10999 1634 11033
rect 1582 10990 1634 10999
rect 1582 10697 1634 10706
rect 1582 10663 1591 10697
rect 1591 10663 1625 10697
rect 1625 10663 1634 10697
rect 1582 10654 1634 10663
rect 1582 10361 1634 10370
rect 1582 10327 1591 10361
rect 1591 10327 1625 10361
rect 1625 10327 1634 10361
rect 1582 10318 1634 10327
rect 1582 10025 1634 10034
rect 1582 9991 1591 10025
rect 1591 9991 1625 10025
rect 1625 9991 1634 10025
rect 1582 9982 1634 9991
rect 1582 9689 1634 9698
rect 1582 9655 1591 9689
rect 1591 9655 1625 9689
rect 1625 9655 1634 9689
rect 1582 9646 1634 9655
rect 1582 9353 1634 9362
rect 1582 9319 1591 9353
rect 1591 9319 1625 9353
rect 1625 9319 1634 9353
rect 1582 9310 1634 9319
rect 1582 9017 1634 9026
rect 1582 8983 1591 9017
rect 1591 8983 1625 9017
rect 1625 8983 1634 9017
rect 1582 8974 1634 8983
rect 1582 8681 1634 8690
rect 1582 8647 1591 8681
rect 1591 8647 1625 8681
rect 1625 8647 1634 8681
rect 1582 8638 1634 8647
rect 1582 8345 1634 8354
rect 1582 8311 1591 8345
rect 1591 8311 1625 8345
rect 1625 8311 1634 8345
rect 1582 8302 1634 8311
rect 1582 8009 1634 8018
rect 1582 7975 1591 8009
rect 1591 7975 1625 8009
rect 1625 7975 1634 8009
rect 1582 7966 1634 7975
rect 1582 7673 1634 7682
rect 1582 7639 1591 7673
rect 1591 7639 1625 7673
rect 1625 7639 1634 7673
rect 1582 7630 1634 7639
rect 1582 7337 1634 7346
rect 1582 7303 1591 7337
rect 1591 7303 1625 7337
rect 1625 7303 1634 7337
rect 1582 7294 1634 7303
rect 1582 7001 1634 7010
rect 1582 6967 1591 7001
rect 1591 6967 1625 7001
rect 1625 6967 1634 7001
rect 1582 6958 1634 6967
rect 66186 17753 66238 17762
rect 66186 17719 66195 17753
rect 66195 17719 66229 17753
rect 66229 17719 66238 17753
rect 66186 17710 66238 17719
rect 66186 17417 66238 17426
rect 66186 17383 66195 17417
rect 66195 17383 66229 17417
rect 66229 17383 66238 17417
rect 66186 17374 66238 17383
rect 66186 17081 66238 17090
rect 66186 17047 66195 17081
rect 66195 17047 66229 17081
rect 66229 17047 66238 17081
rect 66186 17038 66238 17047
rect 66186 16745 66238 16754
rect 66186 16711 66195 16745
rect 66195 16711 66229 16745
rect 66229 16711 66238 16745
rect 66186 16702 66238 16711
rect 66186 16409 66238 16418
rect 66186 16375 66195 16409
rect 66195 16375 66229 16409
rect 66229 16375 66238 16409
rect 66186 16366 66238 16375
rect 66186 16073 66238 16082
rect 66186 16039 66195 16073
rect 66195 16039 66229 16073
rect 66229 16039 66238 16073
rect 66186 16030 66238 16039
rect 66186 15737 66238 15746
rect 66186 15703 66195 15737
rect 66195 15703 66229 15737
rect 66229 15703 66238 15737
rect 66186 15694 66238 15703
rect 66186 15401 66238 15410
rect 66186 15367 66195 15401
rect 66195 15367 66229 15401
rect 66229 15367 66238 15401
rect 66186 15358 66238 15367
rect 66186 15065 66238 15074
rect 66186 15031 66195 15065
rect 66195 15031 66229 15065
rect 66229 15031 66238 15065
rect 66186 15022 66238 15031
rect 66186 14729 66238 14738
rect 66186 14695 66195 14729
rect 66195 14695 66229 14729
rect 66229 14695 66238 14729
rect 66186 14686 66238 14695
rect 66186 14393 66238 14402
rect 66186 14359 66195 14393
rect 66195 14359 66229 14393
rect 66229 14359 66238 14393
rect 66186 14350 66238 14359
rect 56673 13987 56725 14039
rect 66186 14057 66238 14066
rect 66186 14023 66195 14057
rect 66195 14023 66229 14057
rect 66229 14023 66238 14057
rect 66186 14014 66238 14023
rect 66186 13721 66238 13730
rect 66186 13687 66195 13721
rect 66195 13687 66229 13721
rect 66229 13687 66238 13721
rect 66186 13678 66238 13687
rect 66186 13385 66238 13394
rect 66186 13351 66195 13385
rect 66195 13351 66229 13385
rect 66229 13351 66238 13385
rect 66186 13342 66238 13351
rect 66186 13049 66238 13058
rect 66186 13015 66195 13049
rect 66195 13015 66229 13049
rect 66229 13015 66238 13049
rect 66186 13006 66238 13015
rect 66186 12713 66238 12722
rect 66186 12679 66195 12713
rect 66195 12679 66229 12713
rect 66229 12679 66238 12713
rect 66186 12670 66238 12679
rect 56593 12429 56645 12481
rect 66186 12377 66238 12386
rect 66186 12343 66195 12377
rect 66195 12343 66229 12377
rect 66229 12343 66238 12377
rect 66186 12334 66238 12343
rect 66186 12041 66238 12050
rect 66186 12007 66195 12041
rect 66195 12007 66229 12041
rect 66229 12007 66238 12041
rect 66186 11998 66238 12007
rect 66186 11705 66238 11714
rect 66186 11671 66195 11705
rect 66195 11671 66229 11705
rect 66229 11671 66238 11705
rect 66186 11662 66238 11671
rect 66186 11369 66238 11378
rect 66186 11335 66195 11369
rect 66195 11335 66229 11369
rect 66229 11335 66238 11369
rect 66186 11326 66238 11335
rect 56513 11159 56565 11211
rect 66186 11033 66238 11042
rect 66186 10999 66195 11033
rect 66195 10999 66229 11033
rect 66229 10999 66238 11033
rect 66186 10990 66238 10999
rect 66186 10697 66238 10706
rect 66186 10663 66195 10697
rect 66195 10663 66229 10697
rect 66229 10663 66238 10697
rect 66186 10654 66238 10663
rect 66186 10361 66238 10370
rect 66186 10327 66195 10361
rect 66195 10327 66229 10361
rect 66229 10327 66238 10361
rect 66186 10318 66238 10327
rect 66186 10025 66238 10034
rect 66186 9991 66195 10025
rect 66195 9991 66229 10025
rect 66229 9991 66238 10025
rect 66186 9982 66238 9991
rect 56433 9601 56485 9653
rect 66186 9689 66238 9698
rect 66186 9655 66195 9689
rect 66195 9655 66229 9689
rect 66229 9655 66238 9689
rect 66186 9646 66238 9655
rect 66186 9353 66238 9362
rect 66186 9319 66195 9353
rect 66195 9319 66229 9353
rect 66229 9319 66238 9353
rect 66186 9310 66238 9319
rect 66186 9017 66238 9026
rect 66186 8983 66195 9017
rect 66195 8983 66229 9017
rect 66229 8983 66238 9017
rect 66186 8974 66238 8983
rect 66186 8681 66238 8690
rect 66186 8647 66195 8681
rect 66195 8647 66229 8681
rect 66229 8647 66238 8681
rect 66186 8638 66238 8647
rect 56353 8331 56405 8383
rect 66186 8345 66238 8354
rect 66186 8311 66195 8345
rect 66195 8311 66229 8345
rect 66229 8311 66238 8345
rect 66186 8302 66238 8311
rect 66186 8009 66238 8018
rect 66186 7975 66195 8009
rect 66195 7975 66229 8009
rect 66229 7975 66238 8009
rect 66186 7966 66238 7975
rect 66186 7673 66238 7682
rect 66186 7639 66195 7673
rect 66195 7639 66229 7673
rect 66229 7639 66238 7673
rect 66186 7630 66238 7639
rect 66186 7337 66238 7346
rect 66186 7303 66195 7337
rect 66195 7303 66229 7337
rect 66229 7303 66238 7337
rect 66186 7294 66238 7303
rect 66186 7001 66238 7010
rect 66186 6967 66195 7001
rect 66195 6967 66229 7001
rect 66229 6967 66238 7001
rect 66186 6958 66238 6967
rect 56273 6773 56325 6825
rect 1582 6665 1634 6674
rect 1582 6631 1591 6665
rect 1591 6631 1625 6665
rect 1625 6631 1634 6665
rect 1582 6622 1634 6631
rect 66186 6665 66238 6674
rect 66186 6631 66195 6665
rect 66195 6631 66229 6665
rect 66229 6631 66238 6665
rect 66186 6622 66238 6631
rect 1582 6329 1634 6338
rect 1582 6295 1591 6329
rect 1591 6295 1625 6329
rect 1625 6295 1634 6329
rect 1582 6286 1634 6295
rect 66186 6329 66238 6338
rect 66186 6295 66195 6329
rect 66195 6295 66229 6329
rect 66229 6295 66238 6329
rect 66186 6286 66238 6295
rect 1582 5993 1634 6002
rect 1582 5959 1591 5993
rect 1591 5959 1625 5993
rect 1625 5959 1634 5993
rect 1582 5950 1634 5959
rect 66186 5993 66238 6002
rect 66186 5959 66195 5993
rect 66195 5959 66229 5993
rect 66229 5959 66238 5993
rect 66186 5950 66238 5959
rect 1582 5657 1634 5666
rect 1582 5623 1591 5657
rect 1591 5623 1625 5657
rect 1625 5623 1634 5657
rect 1582 5614 1634 5623
rect 66186 5657 66238 5666
rect 66186 5623 66195 5657
rect 66195 5623 66229 5657
rect 66229 5623 66238 5657
rect 66186 5614 66238 5623
rect 1582 5321 1634 5330
rect 1582 5287 1591 5321
rect 1591 5287 1625 5321
rect 1625 5287 1634 5321
rect 1582 5278 1634 5287
rect 66186 5321 66238 5330
rect 66186 5287 66195 5321
rect 66195 5287 66229 5321
rect 66229 5287 66238 5321
rect 66186 5278 66238 5287
rect 1582 4985 1634 4994
rect 1582 4951 1591 4985
rect 1591 4951 1625 4985
rect 1625 4951 1634 4985
rect 1582 4942 1634 4951
rect 66186 4985 66238 4994
rect 66186 4951 66195 4985
rect 66195 4951 66229 4985
rect 66229 4951 66238 4985
rect 66186 4942 66238 4951
rect 1582 4649 1634 4658
rect 1582 4615 1591 4649
rect 1591 4615 1625 4649
rect 1625 4615 1634 4649
rect 1582 4606 1634 4615
rect 66186 4649 66238 4658
rect 66186 4615 66195 4649
rect 66195 4615 66229 4649
rect 66229 4615 66238 4649
rect 66186 4606 66238 4615
rect 1582 4313 1634 4322
rect 1582 4279 1591 4313
rect 1591 4279 1625 4313
rect 1625 4279 1634 4313
rect 1582 4270 1634 4279
rect 66186 4313 66238 4322
rect 66186 4279 66195 4313
rect 66195 4279 66229 4313
rect 66229 4279 66238 4313
rect 66186 4270 66238 4279
rect 1582 3977 1634 3986
rect 1582 3943 1591 3977
rect 1591 3943 1625 3977
rect 1625 3943 1634 3977
rect 1582 3934 1634 3943
rect 66186 3977 66238 3986
rect 66186 3943 66195 3977
rect 66195 3943 66229 3977
rect 66229 3943 66238 3977
rect 66186 3934 66238 3943
rect 1582 3641 1634 3650
rect 1582 3607 1591 3641
rect 1591 3607 1625 3641
rect 1625 3607 1634 3641
rect 1582 3598 1634 3607
rect 66186 3641 66238 3650
rect 66186 3607 66195 3641
rect 66195 3607 66229 3641
rect 66229 3607 66238 3641
rect 66186 3598 66238 3607
rect 1582 3305 1634 3314
rect 1582 3271 1591 3305
rect 1591 3271 1625 3305
rect 1625 3271 1634 3305
rect 1582 3262 1634 3271
rect 66186 3305 66238 3314
rect 66186 3271 66195 3305
rect 66195 3271 66229 3305
rect 66229 3271 66238 3305
rect 66186 3262 66238 3271
rect 1582 2969 1634 2978
rect 1582 2935 1591 2969
rect 1591 2935 1625 2969
rect 1625 2935 1634 2969
rect 1582 2926 1634 2935
rect 66186 2969 66238 2978
rect 66186 2935 66195 2969
rect 66195 2935 66229 2969
rect 66229 2935 66238 2969
rect 66186 2926 66238 2935
rect 1582 2633 1634 2642
rect 1582 2599 1591 2633
rect 1591 2599 1625 2633
rect 1625 2599 1634 2633
rect 1582 2590 1634 2599
rect 66186 2633 66238 2642
rect 66186 2599 66195 2633
rect 66195 2599 66229 2633
rect 66229 2599 66238 2633
rect 66186 2590 66238 2599
rect 1582 2297 1634 2306
rect 1582 2263 1591 2297
rect 1591 2263 1625 2297
rect 1625 2263 1634 2297
rect 1582 2254 1634 2263
rect 66186 2297 66238 2306
rect 66186 2263 66195 2297
rect 66195 2263 66229 2297
rect 66229 2263 66238 2297
rect 66186 2254 66238 2263
rect 1582 1961 1634 1970
rect 1582 1927 1591 1961
rect 1591 1927 1625 1961
rect 1625 1927 1634 1961
rect 1582 1918 1634 1927
rect 66186 1961 66238 1970
rect 66186 1927 66195 1961
rect 66195 1927 66229 1961
rect 66229 1927 66238 1961
rect 66186 1918 66238 1927
rect 1918 1625 1970 1634
rect 3598 1625 3650 1634
rect 5278 1625 5330 1634
rect 6958 1625 7010 1634
rect 8638 1625 8690 1634
rect 10318 1625 10370 1634
rect 11998 1625 12050 1634
rect 13678 1625 13730 1634
rect 15358 1625 15410 1634
rect 17038 1625 17090 1634
rect 18718 1625 18770 1634
rect 20398 1625 20450 1634
rect 22078 1625 22130 1634
rect 23758 1625 23810 1634
rect 25438 1625 25490 1634
rect 27118 1625 27170 1634
rect 28798 1625 28850 1634
rect 30478 1625 30530 1634
rect 32158 1625 32210 1634
rect 33838 1625 33890 1634
rect 35518 1625 35570 1634
rect 37198 1625 37250 1634
rect 38878 1625 38930 1634
rect 40558 1625 40610 1634
rect 42238 1625 42290 1634
rect 43918 1625 43970 1634
rect 45598 1625 45650 1634
rect 47278 1625 47330 1634
rect 48958 1625 49010 1634
rect 50638 1625 50690 1634
rect 52318 1625 52370 1634
rect 53998 1625 54050 1634
rect 55678 1625 55730 1634
rect 57358 1625 57410 1634
rect 59038 1625 59090 1634
rect 60718 1625 60770 1634
rect 62398 1625 62450 1634
rect 64078 1625 64130 1634
rect 65758 1625 65810 1634
rect 1918 1591 1927 1625
rect 1927 1591 1961 1625
rect 1961 1591 1970 1625
rect 3598 1591 3607 1625
rect 3607 1591 3641 1625
rect 3641 1591 3650 1625
rect 5278 1591 5287 1625
rect 5287 1591 5321 1625
rect 5321 1591 5330 1625
rect 6958 1591 6967 1625
rect 6967 1591 7001 1625
rect 7001 1591 7010 1625
rect 8638 1591 8647 1625
rect 8647 1591 8681 1625
rect 8681 1591 8690 1625
rect 10318 1591 10327 1625
rect 10327 1591 10361 1625
rect 10361 1591 10370 1625
rect 11998 1591 12007 1625
rect 12007 1591 12041 1625
rect 12041 1591 12050 1625
rect 13678 1591 13687 1625
rect 13687 1591 13721 1625
rect 13721 1591 13730 1625
rect 15358 1591 15367 1625
rect 15367 1591 15401 1625
rect 15401 1591 15410 1625
rect 17038 1591 17047 1625
rect 17047 1591 17081 1625
rect 17081 1591 17090 1625
rect 18718 1591 18727 1625
rect 18727 1591 18761 1625
rect 18761 1591 18770 1625
rect 20398 1591 20407 1625
rect 20407 1591 20441 1625
rect 20441 1591 20450 1625
rect 22078 1591 22087 1625
rect 22087 1591 22121 1625
rect 22121 1591 22130 1625
rect 23758 1591 23767 1625
rect 23767 1591 23801 1625
rect 23801 1591 23810 1625
rect 25438 1591 25447 1625
rect 25447 1591 25481 1625
rect 25481 1591 25490 1625
rect 27118 1591 27127 1625
rect 27127 1591 27161 1625
rect 27161 1591 27170 1625
rect 28798 1591 28807 1625
rect 28807 1591 28841 1625
rect 28841 1591 28850 1625
rect 30478 1591 30487 1625
rect 30487 1591 30521 1625
rect 30521 1591 30530 1625
rect 32158 1591 32167 1625
rect 32167 1591 32201 1625
rect 32201 1591 32210 1625
rect 33838 1591 33847 1625
rect 33847 1591 33881 1625
rect 33881 1591 33890 1625
rect 35518 1591 35527 1625
rect 35527 1591 35561 1625
rect 35561 1591 35570 1625
rect 37198 1591 37207 1625
rect 37207 1591 37241 1625
rect 37241 1591 37250 1625
rect 38878 1591 38887 1625
rect 38887 1591 38921 1625
rect 38921 1591 38930 1625
rect 40558 1591 40567 1625
rect 40567 1591 40601 1625
rect 40601 1591 40610 1625
rect 42238 1591 42247 1625
rect 42247 1591 42281 1625
rect 42281 1591 42290 1625
rect 43918 1591 43927 1625
rect 43927 1591 43961 1625
rect 43961 1591 43970 1625
rect 45598 1591 45607 1625
rect 45607 1591 45641 1625
rect 45641 1591 45650 1625
rect 47278 1591 47287 1625
rect 47287 1591 47321 1625
rect 47321 1591 47330 1625
rect 48958 1591 48967 1625
rect 48967 1591 49001 1625
rect 49001 1591 49010 1625
rect 50638 1591 50647 1625
rect 50647 1591 50681 1625
rect 50681 1591 50690 1625
rect 52318 1591 52327 1625
rect 52327 1591 52361 1625
rect 52361 1591 52370 1625
rect 53998 1591 54007 1625
rect 54007 1591 54041 1625
rect 54041 1591 54050 1625
rect 55678 1591 55687 1625
rect 55687 1591 55721 1625
rect 55721 1591 55730 1625
rect 57358 1591 57367 1625
rect 57367 1591 57401 1625
rect 57401 1591 57410 1625
rect 59038 1591 59047 1625
rect 59047 1591 59081 1625
rect 59081 1591 59090 1625
rect 60718 1591 60727 1625
rect 60727 1591 60761 1625
rect 60761 1591 60770 1625
rect 62398 1591 62407 1625
rect 62407 1591 62441 1625
rect 62441 1591 62450 1625
rect 64078 1591 64087 1625
rect 64087 1591 64121 1625
rect 64121 1591 64130 1625
rect 65758 1591 65767 1625
rect 65767 1591 65801 1625
rect 65801 1591 65810 1625
rect 1918 1582 1970 1591
rect 3598 1582 3650 1591
rect 5278 1582 5330 1591
rect 6958 1582 7010 1591
rect 8638 1582 8690 1591
rect 10318 1582 10370 1591
rect 11998 1582 12050 1591
rect 13678 1582 13730 1591
rect 15358 1582 15410 1591
rect 17038 1582 17090 1591
rect 18718 1582 18770 1591
rect 20398 1582 20450 1591
rect 22078 1582 22130 1591
rect 23758 1582 23810 1591
rect 25438 1582 25490 1591
rect 27118 1582 27170 1591
rect 28798 1582 28850 1591
rect 30478 1582 30530 1591
rect 32158 1582 32210 1591
rect 33838 1582 33890 1591
rect 35518 1582 35570 1591
rect 37198 1582 37250 1591
rect 38878 1582 38930 1591
rect 40558 1582 40610 1591
rect 42238 1582 42290 1591
rect 43918 1582 43970 1591
rect 45598 1582 45650 1591
rect 47278 1582 47330 1591
rect 48958 1582 49010 1591
rect 50638 1582 50690 1591
rect 52318 1582 52370 1591
rect 53998 1582 54050 1591
rect 55678 1582 55730 1591
rect 57358 1582 57410 1591
rect 59038 1582 59090 1591
rect 60718 1582 60770 1591
rect 62398 1582 62450 1591
rect 64078 1582 64130 1591
rect 65758 1582 65810 1591
<< metal2 >>
rect 1496 50692 1720 51242
rect 1916 51158 1972 51167
rect 1916 51093 1972 51102
rect 3596 51158 3652 51167
rect 3596 51093 3652 51102
rect 5276 51158 5332 51167
rect 5276 51093 5332 51102
rect 6956 51158 7012 51167
rect 6956 51093 7012 51102
rect 8636 51158 8692 51167
rect 8636 51093 8692 51102
rect 10316 51158 10372 51167
rect 10316 51093 10372 51102
rect 11996 51158 12052 51167
rect 11996 51093 12052 51102
rect 13676 51158 13732 51167
rect 13676 51093 13732 51102
rect 15356 51158 15412 51167
rect 15356 51093 15412 51102
rect 17036 51158 17092 51167
rect 17036 51093 17092 51102
rect 18716 51158 18772 51167
rect 18716 51093 18772 51102
rect 20396 51158 20452 51167
rect 20396 51093 20452 51102
rect 22076 51158 22132 51167
rect 22076 51093 22132 51102
rect 23756 51158 23812 51167
rect 23756 51093 23812 51102
rect 25436 51158 25492 51167
rect 25436 51093 25492 51102
rect 27116 51158 27172 51167
rect 27116 51093 27172 51102
rect 28796 51158 28852 51167
rect 28796 51093 28852 51102
rect 30476 51158 30532 51167
rect 30476 51093 30532 51102
rect 32156 51158 32212 51167
rect 32156 51093 32212 51102
rect 33836 51158 33892 51167
rect 33836 51093 33892 51102
rect 35516 51158 35572 51167
rect 35516 51093 35572 51102
rect 37196 51158 37252 51167
rect 37196 51093 37252 51102
rect 38876 51158 38932 51167
rect 38876 51093 38932 51102
rect 40556 51158 40612 51167
rect 40556 51093 40612 51102
rect 42236 51158 42292 51167
rect 42236 51093 42292 51102
rect 43916 51158 43972 51167
rect 43916 51093 43972 51102
rect 45596 51158 45652 51167
rect 45596 51093 45652 51102
rect 47276 51158 47332 51167
rect 47276 51093 47332 51102
rect 48956 51158 49012 51167
rect 48956 51093 49012 51102
rect 50636 51158 50692 51167
rect 50636 51093 50692 51102
rect 52316 51158 52372 51167
rect 52316 51093 52372 51102
rect 53996 51158 54052 51167
rect 53996 51093 54052 51102
rect 55676 51158 55732 51167
rect 55676 51093 55732 51102
rect 57356 51158 57412 51167
rect 57356 51093 57412 51102
rect 59036 51158 59092 51167
rect 59036 51093 59092 51102
rect 60716 51158 60772 51167
rect 60716 51093 60772 51102
rect 62396 51158 62452 51167
rect 62396 51093 62452 51102
rect 64076 51158 64132 51167
rect 64076 51093 64132 51102
rect 65756 51158 65812 51167
rect 65756 51093 65812 51102
rect 1496 50636 1580 50692
rect 1636 50636 1720 50692
rect 1496 50354 1720 50636
rect 1496 50302 1582 50354
rect 1634 50302 1720 50354
rect 1496 50018 1720 50302
rect 66100 50692 66324 51242
rect 66100 50636 66184 50692
rect 66240 50636 66324 50692
rect 66100 50354 66324 50636
rect 66100 50302 66186 50354
rect 66238 50302 66324 50354
rect 1496 49966 1582 50018
rect 1634 49966 1720 50018
rect 1496 49682 1720 49966
rect 56872 50010 56928 50019
rect 56872 49945 56928 49954
rect 66100 50018 66324 50302
rect 66100 49966 66186 50018
rect 66238 49966 66324 50018
rect 53282 49754 53338 49763
rect 53282 49689 53338 49698
rect 54450 49754 54506 49763
rect 54450 49689 54506 49698
rect 1496 49630 1582 49682
rect 1634 49630 1720 49682
rect 1496 49346 1720 49630
rect 1496 49294 1582 49346
rect 1634 49294 1720 49346
rect 1496 49012 1720 49294
rect 1496 48956 1580 49012
rect 1636 48956 1720 49012
rect 1496 48674 1720 48956
rect 1496 48622 1582 48674
rect 1634 48622 1720 48674
rect 1496 48338 1720 48622
rect 1496 48286 1582 48338
rect 1634 48286 1720 48338
rect 1496 48002 1720 48286
rect 1496 47950 1582 48002
rect 1634 47950 1720 48002
rect 1496 47666 1720 47950
rect 1496 47614 1582 47666
rect 1634 47614 1720 47666
rect 1496 47332 1720 47614
rect 1496 47276 1580 47332
rect 1636 47276 1720 47332
rect 1496 46994 1720 47276
rect 1496 46942 1582 46994
rect 1634 46942 1720 46994
rect 1496 46658 1720 46942
rect 56886 48633 56914 49945
rect 66100 49682 66324 49966
rect 66100 49630 66186 49682
rect 66238 49630 66324 49682
rect 66100 49346 66324 49630
rect 66100 49294 66186 49346
rect 66238 49294 66324 49346
rect 66100 49012 66324 49294
rect 66100 48956 66184 49012
rect 66240 48956 66324 49012
rect 65056 48790 65112 48799
rect 65056 48725 65112 48734
rect 61759 48685 61815 48694
rect 56886 48605 56984 48633
rect 61759 48620 61815 48629
rect 66100 48674 66324 48956
rect 66100 48622 66186 48674
rect 66238 48622 66324 48674
rect 23983 46889 24039 46898
rect 23983 46824 24039 46833
rect 26479 46889 26535 46898
rect 26479 46824 26535 46833
rect 28975 46889 29031 46898
rect 28975 46824 29031 46833
rect 31471 46889 31527 46898
rect 31471 46824 31527 46833
rect 33967 46889 34023 46898
rect 33967 46824 34023 46833
rect 36463 46889 36519 46898
rect 36463 46824 36519 46833
rect 38959 46889 39015 46898
rect 38959 46824 39015 46833
rect 41455 46889 41511 46898
rect 41455 46824 41511 46833
rect 1496 46606 1582 46658
rect 1634 46606 1720 46658
rect 1496 46322 1720 46606
rect 1496 46270 1582 46322
rect 1634 46270 1720 46322
rect 1496 45986 1720 46270
rect 1496 45934 1582 45986
rect 1634 45934 1720 45986
rect 1496 45652 1720 45934
rect 1496 45596 1580 45652
rect 1636 45596 1720 45652
rect 1496 45314 1720 45596
rect 1496 45262 1582 45314
rect 1634 45262 1720 45314
rect 1496 44978 1720 45262
rect 1496 44926 1582 44978
rect 1634 44926 1720 44978
rect 1496 44642 1720 44926
rect 1496 44590 1582 44642
rect 1634 44590 1720 44642
rect 1496 44306 1720 44590
rect 46067 44389 46123 44398
rect 46067 44324 46123 44333
rect 1496 44254 1582 44306
rect 1634 44254 1720 44306
rect 1496 43972 1720 44254
rect 1496 43916 1580 43972
rect 1636 43916 1720 43972
rect 1496 43634 1720 43916
rect 1496 43582 1582 43634
rect 1634 43582 1720 43634
rect 1496 43298 1720 43582
rect 1496 43246 1582 43298
rect 1634 43246 1720 43298
rect 1496 42962 1720 43246
rect 1496 42910 1582 42962
rect 1634 42910 1720 42962
rect 1496 42626 1720 42910
rect 1496 42574 1582 42626
rect 1634 42574 1720 42626
rect 1496 42292 1720 42574
rect 1496 42236 1580 42292
rect 1636 42236 1720 42292
rect 1496 41954 1720 42236
rect 1496 41902 1582 41954
rect 1634 41902 1720 41954
rect 1496 41618 1720 41902
rect 1496 41566 1582 41618
rect 1634 41566 1720 41618
rect 1496 41282 1720 41566
rect 1496 41230 1582 41282
rect 1634 41230 1720 41282
rect 1496 40946 1720 41230
rect 1496 40894 1582 40946
rect 1634 40894 1720 40946
rect 1496 40612 1720 40894
rect 46081 40704 46109 44324
rect 46191 42991 46247 43000
rect 46191 42926 46247 42935
rect 46205 40704 46233 42926
rect 49252 41577 49308 41586
rect 49252 41512 49308 41521
rect 1496 40556 1580 40612
rect 1636 40556 1720 40612
rect 1496 40274 1720 40556
rect 1496 40222 1582 40274
rect 1634 40222 1720 40274
rect 49266 40227 49294 41512
rect 1496 39938 1720 40222
rect 46769 40153 46825 40162
rect 46769 40088 46825 40097
rect 48660 40141 48716 40150
rect 48660 40076 48716 40085
rect 1496 39886 1582 39938
rect 1634 39886 1720 39938
rect 1496 39602 1720 39886
rect 1496 39550 1582 39602
rect 1634 39550 1720 39602
rect 1496 39266 1720 39550
rect 1496 39214 1582 39266
rect 1634 39214 1720 39266
rect 1496 38932 1720 39214
rect 1496 38876 1580 38932
rect 1636 38876 1720 38932
rect 1496 38594 1720 38876
rect 1496 38542 1582 38594
rect 1634 38542 1720 38594
rect 1496 38258 1720 38542
rect 1496 38206 1582 38258
rect 1634 38206 1720 38258
rect 1496 37922 1720 38206
rect 1496 37870 1582 37922
rect 1634 37870 1720 37922
rect 1496 37586 1720 37870
rect 1496 37534 1582 37586
rect 1634 37534 1720 37586
rect 1496 37252 1720 37534
rect 1496 37196 1580 37252
rect 1636 37196 1720 37252
rect 1496 36914 1720 37196
rect 1496 36862 1582 36914
rect 1634 36862 1720 36914
rect 1496 36578 1720 36862
rect 1496 36526 1582 36578
rect 1634 36526 1720 36578
rect 1496 36242 1720 36526
rect 1496 36190 1582 36242
rect 1634 36190 1720 36242
rect 1496 35906 1720 36190
rect 1496 35854 1582 35906
rect 1634 35854 1720 35906
rect 1496 35572 1720 35854
rect 1496 35516 1580 35572
rect 1636 35516 1720 35572
rect 1496 35234 1720 35516
rect 1496 35182 1582 35234
rect 1634 35182 1720 35234
rect 1496 34898 1720 35182
rect 1496 34846 1582 34898
rect 1634 34846 1720 34898
rect 1496 34562 1720 34846
rect 1496 34510 1582 34562
rect 1634 34510 1720 34562
rect 1496 34226 1720 34510
rect 1496 34174 1582 34226
rect 1634 34174 1720 34226
rect 1496 33892 1720 34174
rect 1496 33836 1580 33892
rect 1636 33836 1720 33892
rect 1496 33554 1720 33836
rect 1496 33502 1582 33554
rect 1634 33502 1720 33554
rect 1496 33218 1720 33502
rect 1496 33166 1582 33218
rect 1634 33166 1720 33218
rect 1496 32882 1720 33166
rect 1496 32830 1582 32882
rect 1634 32830 1720 32882
rect 1496 32546 1720 32830
rect 1496 32494 1582 32546
rect 1634 32494 1720 32546
rect 1496 32212 1720 32494
rect 1496 32156 1580 32212
rect 1636 32156 1720 32212
rect 1496 31874 1720 32156
rect 1496 31822 1582 31874
rect 1634 31822 1720 31874
rect 1496 31538 1720 31822
rect 1496 31486 1582 31538
rect 1634 31486 1720 31538
rect 1496 31202 1720 31486
rect 1496 31150 1582 31202
rect 1634 31150 1720 31202
rect 1496 30866 1720 31150
rect 1496 30814 1582 30866
rect 1634 30814 1720 30866
rect 1496 30532 1720 30814
rect 1496 30476 1580 30532
rect 1636 30476 1720 30532
rect 1496 30194 1720 30476
rect 9810 30276 9866 30285
rect 9810 30211 9866 30220
rect 1496 30142 1582 30194
rect 1634 30142 1720 30194
rect 1496 29858 1720 30142
rect 10755 30205 10811 30214
rect 10755 30140 10811 30149
rect 11409 30205 11465 30214
rect 11409 30140 11465 30149
rect 1496 29806 1582 29858
rect 1634 29806 1720 29858
rect 1496 29522 1720 29806
rect 1496 29470 1582 29522
rect 1634 29470 1720 29522
rect 1496 29186 1720 29470
rect 1496 29134 1582 29186
rect 1634 29134 1720 29186
rect 1496 28852 1720 29134
rect 1496 28796 1580 28852
rect 1636 28796 1720 28852
rect 1496 28514 1720 28796
rect 10755 28647 10811 28656
rect 1496 28462 1582 28514
rect 1634 28462 1720 28514
rect 9810 28576 9866 28585
rect 10755 28582 10811 28591
rect 11329 28647 11385 28656
rect 11329 28582 11385 28591
rect 9810 28511 9866 28520
rect 1496 28178 1720 28462
rect 1496 28126 1582 28178
rect 1634 28126 1720 28178
rect 1496 27842 1720 28126
rect 1496 27790 1582 27842
rect 1634 27790 1720 27842
rect 1496 27506 1720 27790
rect 1496 27454 1582 27506
rect 1634 27454 1720 27506
rect 1496 27172 1720 27454
rect 9810 27448 9866 27457
rect 9810 27383 9866 27392
rect 10755 27377 10811 27386
rect 10755 27312 10811 27321
rect 11249 27377 11305 27386
rect 11249 27312 11305 27321
rect 1496 27116 1580 27172
rect 1636 27116 1720 27172
rect 1496 26834 1720 27116
rect 1496 26782 1582 26834
rect 1634 26782 1720 26834
rect 1496 26498 1720 26782
rect 1496 26446 1582 26498
rect 1634 26446 1720 26498
rect 1496 26162 1720 26446
rect 1496 26110 1582 26162
rect 1634 26110 1720 26162
rect 1496 25826 1720 26110
rect 1496 25774 1582 25826
rect 1634 25774 1720 25826
rect 1496 25492 1720 25774
rect 10755 25819 10811 25828
rect 9810 25748 9866 25757
rect 10755 25754 10811 25763
rect 11169 25819 11225 25828
rect 11169 25754 11225 25763
rect 9810 25683 9866 25692
rect 1496 25436 1580 25492
rect 1636 25436 1720 25492
rect 1496 25154 1720 25436
rect 1496 25102 1582 25154
rect 1634 25102 1720 25154
rect 1496 24818 1720 25102
rect 1496 24766 1582 24818
rect 1634 24766 1720 24818
rect 1496 24482 1720 24766
rect 9810 24620 9866 24629
rect 9810 24555 9866 24564
rect 10755 24549 10811 24558
rect 10755 24484 10811 24493
rect 11089 24549 11145 24558
rect 11089 24484 11145 24493
rect 1496 24430 1582 24482
rect 1634 24430 1720 24482
rect 1496 24146 1720 24430
rect 1496 24094 1582 24146
rect 1634 24094 1720 24146
rect 1496 23812 1720 24094
rect 1496 23756 1580 23812
rect 1636 23756 1720 23812
rect 1496 23474 1720 23756
rect 1496 23422 1582 23474
rect 1634 23422 1720 23474
rect 1496 23138 1720 23422
rect 1496 23086 1582 23138
rect 1634 23086 1720 23138
rect 1496 22802 1720 23086
rect 10755 22991 10811 23000
rect 9810 22920 9866 22929
rect 10755 22926 10811 22935
rect 11009 22991 11065 23000
rect 11009 22926 11065 22935
rect 9810 22855 9866 22864
rect 1496 22750 1582 22802
rect 1634 22750 1720 22802
rect 1496 22466 1720 22750
rect 10892 22664 10948 22673
rect 10892 22599 10948 22608
rect 1496 22414 1582 22466
rect 1634 22414 1720 22466
rect 1496 22132 1720 22414
rect 1496 22076 1580 22132
rect 1636 22076 1720 22132
rect 1496 21794 1720 22076
rect 1496 21742 1582 21794
rect 1634 21742 1720 21794
rect 1496 21458 1720 21742
rect 2495 21527 2551 21536
rect 2495 21462 2551 21471
rect 1496 21406 1582 21458
rect 1634 21406 1720 21458
rect 1496 21122 1720 21406
rect 1496 21070 1582 21122
rect 1634 21070 1720 21122
rect 1496 20786 1720 21070
rect 1496 20734 1582 20786
rect 1634 20734 1720 20786
rect 1496 20452 1720 20734
rect 1496 20396 1580 20452
rect 1636 20396 1720 20452
rect 1496 20114 1720 20396
rect 1496 20062 1582 20114
rect 1634 20062 1720 20114
rect 1496 19778 1720 20062
rect 1496 19726 1582 19778
rect 1634 19726 1720 19778
rect 1496 19442 1720 19726
rect 1496 19390 1582 19442
rect 1634 19390 1720 19442
rect 1496 19106 1720 19390
rect 1496 19054 1582 19106
rect 1634 19054 1720 19106
rect 1496 18772 1720 19054
rect 1496 18716 1580 18772
rect 1636 18716 1720 18772
rect 1496 18434 1720 18716
rect 1496 18382 1582 18434
rect 1634 18382 1720 18434
rect 1496 18098 1720 18382
rect 1496 18046 1582 18098
rect 1634 18046 1720 18098
rect 1496 17762 1720 18046
rect 1496 17710 1582 17762
rect 1634 17710 1720 17762
rect 1496 17426 1720 17710
rect 1496 17374 1582 17426
rect 1634 17374 1720 17426
rect 1496 17092 1720 17374
rect 1496 17036 1580 17092
rect 1636 17036 1720 17092
rect 1496 16754 1720 17036
rect 1496 16702 1582 16754
rect 1634 16702 1720 16754
rect 1496 16418 1720 16702
rect 1496 16366 1582 16418
rect 1634 16366 1720 16418
rect 1496 16082 1720 16366
rect 1496 16030 1582 16082
rect 1634 16030 1720 16082
rect 1496 15746 1720 16030
rect 1496 15694 1582 15746
rect 1634 15694 1720 15746
rect 1496 15412 1720 15694
rect 1496 15356 1580 15412
rect 1636 15356 1720 15412
rect 1496 15074 1720 15356
rect 1496 15022 1582 15074
rect 1634 15022 1720 15074
rect 1496 14738 1720 15022
rect 1496 14686 1582 14738
rect 1634 14686 1720 14738
rect 1496 14402 1720 14686
rect 1496 14350 1582 14402
rect 1634 14350 1720 14402
rect 1496 14066 1720 14350
rect 1496 14014 1582 14066
rect 1634 14014 1720 14066
rect 1496 13732 1720 14014
rect 1496 13676 1580 13732
rect 1636 13676 1720 13732
rect 1496 13394 1720 13676
rect 1496 13342 1582 13394
rect 1634 13342 1720 13394
rect 1496 13058 1720 13342
rect 1496 13006 1582 13058
rect 1634 13006 1720 13058
rect 1496 12722 1720 13006
rect 10808 13005 10864 13014
rect 10808 12940 10864 12949
rect 1496 12670 1582 12722
rect 1634 12670 1720 12722
rect 1496 12386 1720 12670
rect 1496 12334 1582 12386
rect 1634 12334 1720 12386
rect 1496 12052 1720 12334
rect 1496 11996 1580 12052
rect 1636 11996 1720 12052
rect 1496 11714 1720 11996
rect 1496 11662 1582 11714
rect 1634 11662 1720 11714
rect 1496 11378 1720 11662
rect 1496 11326 1582 11378
rect 1634 11326 1720 11378
rect 1496 11042 1720 11326
rect 1496 10990 1582 11042
rect 1634 10990 1720 11042
rect 1496 10706 1720 10990
rect 1496 10654 1582 10706
rect 1634 10654 1720 10706
rect 1496 10372 1720 10654
rect 1496 10316 1580 10372
rect 1636 10316 1720 10372
rect 1496 10034 1720 10316
rect 10808 10177 10864 10186
rect 10808 10112 10864 10121
rect 1496 9982 1582 10034
rect 1634 9982 1720 10034
rect 1496 9698 1720 9982
rect 1496 9646 1582 9698
rect 1634 9646 1720 9698
rect 1496 9362 1720 9646
rect 1496 9310 1582 9362
rect 1634 9310 1720 9362
rect 1496 9026 1720 9310
rect 1496 8974 1582 9026
rect 1634 8974 1720 9026
rect 1496 8692 1720 8974
rect 10808 8763 10864 8772
rect 10808 8698 10864 8707
rect 1496 8636 1580 8692
rect 1636 8636 1720 8692
rect 1496 8354 1720 8636
rect 1496 8302 1582 8354
rect 1634 8302 1720 8354
rect 1496 8018 1720 8302
rect 1496 7966 1582 8018
rect 1634 7966 1720 8018
rect 1496 7682 1720 7966
rect 1496 7630 1582 7682
rect 1634 7630 1720 7682
rect 1496 7346 1720 7630
rect 1496 7294 1582 7346
rect 1634 7294 1720 7346
rect 1496 7012 1720 7294
rect 1496 6956 1580 7012
rect 1636 6956 1720 7012
rect 1496 6674 1720 6956
rect 1496 6622 1582 6674
rect 1634 6622 1720 6674
rect 1496 6338 1720 6622
rect 1496 6286 1582 6338
rect 1634 6286 1720 6338
rect 1496 6002 1720 6286
rect 1496 5950 1582 6002
rect 1634 5950 1720 6002
rect 1496 5666 1720 5950
rect 1496 5614 1582 5666
rect 1634 5614 1720 5666
rect 1496 5332 1720 5614
rect 1496 5276 1580 5332
rect 1636 5276 1720 5332
rect 1496 4994 1720 5276
rect 1496 4942 1582 4994
rect 1634 4942 1720 4994
rect 1496 4658 1720 4942
rect 1496 4606 1582 4658
rect 1634 4606 1720 4658
rect 1496 4322 1720 4606
rect 10906 4507 10934 22599
rect 19020 14491 19076 14500
rect 19020 14426 19076 14435
rect 20911 14479 20967 14488
rect 20911 14414 20967 14423
rect 56886 14377 56914 48605
rect 66100 48338 66324 48622
rect 66100 48286 66186 48338
rect 66238 48286 66324 48338
rect 66100 48002 66324 48286
rect 66100 47950 66186 48002
rect 66238 47950 66324 48002
rect 66100 47666 66324 47950
rect 66100 47614 66186 47666
rect 66238 47614 66324 47666
rect 66100 47332 66324 47614
rect 66100 47276 66184 47332
rect 66240 47276 66324 47332
rect 66100 46994 66324 47276
rect 66100 46942 66186 46994
rect 66238 46942 66324 46994
rect 66100 46658 66324 46942
rect 66100 46606 66186 46658
rect 66238 46606 66324 46658
rect 66100 46322 66324 46606
rect 66100 46270 66186 46322
rect 66238 46270 66324 46322
rect 66100 45986 66324 46270
rect 66100 45934 66186 45986
rect 66238 45934 66324 45986
rect 66100 45652 66324 45934
rect 66100 45596 66184 45652
rect 66240 45596 66324 45652
rect 66100 45314 66324 45596
rect 66100 45262 66186 45314
rect 66238 45262 66324 45314
rect 66100 44978 66324 45262
rect 66100 44926 66186 44978
rect 66238 44926 66324 44978
rect 66100 44642 66324 44926
rect 66100 44590 66186 44642
rect 66238 44590 66324 44642
rect 56956 44389 57012 44398
rect 56956 44324 57012 44333
rect 66100 44306 66324 44590
rect 66100 44254 66186 44306
rect 66238 44254 66324 44306
rect 66100 43972 66324 44254
rect 66100 43916 66184 43972
rect 66240 43916 66324 43972
rect 66100 43634 66324 43916
rect 66100 43582 66186 43634
rect 66238 43582 66324 43634
rect 66100 43298 66324 43582
rect 66100 43246 66186 43298
rect 66238 43246 66324 43298
rect 56956 42991 57012 43000
rect 56956 42926 57012 42935
rect 66100 42962 66324 43246
rect 66100 42910 66186 42962
rect 66238 42910 66324 42962
rect 66100 42626 66324 42910
rect 66100 42574 66186 42626
rect 66238 42574 66324 42626
rect 66100 42292 66324 42574
rect 66100 42236 66184 42292
rect 66240 42236 66324 42292
rect 66100 41954 66324 42236
rect 66100 41902 66186 41954
rect 66238 41902 66324 41954
rect 66100 41618 66324 41902
rect 56956 41577 57012 41586
rect 56956 41512 57012 41521
rect 66100 41566 66186 41618
rect 66238 41566 66324 41618
rect 66100 41282 66324 41566
rect 66100 41230 66186 41282
rect 66238 41230 66324 41282
rect 66100 40946 66324 41230
rect 66100 40894 66186 40946
rect 66238 40894 66324 40946
rect 66100 40612 66324 40894
rect 66100 40556 66184 40612
rect 66240 40556 66324 40612
rect 66100 40274 66324 40556
rect 66100 40222 66186 40274
rect 66238 40222 66324 40274
rect 66100 39938 66324 40222
rect 66100 39886 66186 39938
rect 66238 39886 66324 39938
rect 66100 39602 66324 39886
rect 66100 39550 66186 39602
rect 66238 39550 66324 39602
rect 66100 39266 66324 39550
rect 66100 39214 66186 39266
rect 66238 39214 66324 39266
rect 66100 38932 66324 39214
rect 66100 38876 66184 38932
rect 66240 38876 66324 38932
rect 66100 38594 66324 38876
rect 66100 38542 66186 38594
rect 66238 38542 66324 38594
rect 66100 38258 66324 38542
rect 66100 38206 66186 38258
rect 66238 38206 66324 38258
rect 66100 37922 66324 38206
rect 66100 37870 66186 37922
rect 66238 37870 66324 37922
rect 66100 37586 66324 37870
rect 66100 37534 66186 37586
rect 66238 37534 66324 37586
rect 66100 37252 66324 37534
rect 66100 37196 66184 37252
rect 66240 37196 66324 37252
rect 66100 36914 66324 37196
rect 66100 36862 66186 36914
rect 66238 36862 66324 36914
rect 66100 36578 66324 36862
rect 66100 36526 66186 36578
rect 66238 36526 66324 36578
rect 66100 36242 66324 36526
rect 66100 36190 66186 36242
rect 66238 36190 66324 36242
rect 66100 35906 66324 36190
rect 66100 35854 66186 35906
rect 66238 35854 66324 35906
rect 66100 35572 66324 35854
rect 66100 35516 66184 35572
rect 66240 35516 66324 35572
rect 66100 35234 66324 35516
rect 66100 35182 66186 35234
rect 66238 35182 66324 35234
rect 66100 34898 66324 35182
rect 66100 34846 66186 34898
rect 66238 34846 66324 34898
rect 66100 34562 66324 34846
rect 66100 34510 66186 34562
rect 66238 34510 66324 34562
rect 66100 34226 66324 34510
rect 66100 34174 66186 34226
rect 66238 34174 66324 34226
rect 66100 33892 66324 34174
rect 66100 33836 66184 33892
rect 66240 33836 66324 33892
rect 66100 33554 66324 33836
rect 66100 33502 66186 33554
rect 66238 33502 66324 33554
rect 66100 33218 66324 33502
rect 66100 33166 66186 33218
rect 66238 33166 66324 33218
rect 66100 32882 66324 33166
rect 66100 32830 66186 32882
rect 66238 32830 66324 32882
rect 66100 32546 66324 32830
rect 66100 32494 66186 32546
rect 66238 32494 66324 32546
rect 66100 32212 66324 32494
rect 66100 32156 66184 32212
rect 66240 32156 66324 32212
rect 66100 31874 66324 32156
rect 66100 31822 66186 31874
rect 66238 31822 66324 31874
rect 65269 31641 65325 31650
rect 65269 31576 65325 31585
rect 66100 31538 66324 31822
rect 66100 31486 66186 31538
rect 66238 31486 66324 31538
rect 66100 31202 66324 31486
rect 66100 31150 66186 31202
rect 66238 31150 66324 31202
rect 66100 30866 66324 31150
rect 66100 30814 66186 30866
rect 66238 30814 66324 30866
rect 66100 30532 66324 30814
rect 66100 30476 66184 30532
rect 66240 30476 66324 30532
rect 66100 30194 66324 30476
rect 66100 30142 66186 30194
rect 66238 30142 66324 30194
rect 66100 29858 66324 30142
rect 66100 29806 66186 29858
rect 66238 29806 66324 29858
rect 66100 29522 66324 29806
rect 66100 29470 66186 29522
rect 66238 29470 66324 29522
rect 66100 29186 66324 29470
rect 66100 29134 66186 29186
rect 66238 29134 66324 29186
rect 66100 28852 66324 29134
rect 66100 28796 66184 28852
rect 66240 28796 66324 28852
rect 66100 28514 66324 28796
rect 66100 28462 66186 28514
rect 66238 28462 66324 28514
rect 66100 28178 66324 28462
rect 66100 28126 66186 28178
rect 66238 28126 66324 28178
rect 66100 27842 66324 28126
rect 66100 27790 66186 27842
rect 66238 27790 66324 27842
rect 66100 27506 66324 27790
rect 66100 27454 66186 27506
rect 66238 27454 66324 27506
rect 66100 27172 66324 27454
rect 66100 27116 66184 27172
rect 66240 27116 66324 27172
rect 66100 26834 66324 27116
rect 66100 26782 66186 26834
rect 66238 26782 66324 26834
rect 66100 26498 66324 26782
rect 66100 26446 66186 26498
rect 66238 26446 66324 26498
rect 66100 26162 66324 26446
rect 66100 26110 66186 26162
rect 66238 26110 66324 26162
rect 66100 25826 66324 26110
rect 66100 25774 66186 25826
rect 66238 25774 66324 25826
rect 66100 25492 66324 25774
rect 66100 25436 66184 25492
rect 66240 25436 66324 25492
rect 66100 25154 66324 25436
rect 66100 25102 66186 25154
rect 66238 25102 66324 25154
rect 66100 24818 66324 25102
rect 66100 24766 66186 24818
rect 66238 24766 66324 24818
rect 66100 24482 66324 24766
rect 66100 24430 66186 24482
rect 66238 24430 66324 24482
rect 66100 24146 66324 24430
rect 66100 24094 66186 24146
rect 66238 24094 66324 24146
rect 66100 23812 66324 24094
rect 66100 23756 66184 23812
rect 66240 23756 66324 23812
rect 66100 23474 66324 23756
rect 66100 23422 66186 23474
rect 66238 23422 66324 23474
rect 66100 23138 66324 23422
rect 66100 23086 66186 23138
rect 66238 23086 66324 23138
rect 66100 22802 66324 23086
rect 66100 22750 66186 22802
rect 66238 22750 66324 22802
rect 66100 22466 66324 22750
rect 66100 22414 66186 22466
rect 66238 22414 66324 22466
rect 66100 22132 66324 22414
rect 66100 22076 66184 22132
rect 66240 22076 66324 22132
rect 66100 21794 66324 22076
rect 66100 21742 66186 21794
rect 66238 21742 66324 21794
rect 66100 21458 66324 21742
rect 66100 21406 66186 21458
rect 66238 21406 66324 21458
rect 66100 21122 66324 21406
rect 66100 21070 66186 21122
rect 66238 21070 66324 21122
rect 66100 20786 66324 21070
rect 66100 20734 66186 20786
rect 66238 20734 66324 20786
rect 66100 20452 66324 20734
rect 66100 20396 66184 20452
rect 66240 20396 66324 20452
rect 66100 20114 66324 20396
rect 66100 20062 66186 20114
rect 66238 20062 66324 20114
rect 66100 19778 66324 20062
rect 66100 19726 66186 19778
rect 66238 19726 66324 19778
rect 66100 19442 66324 19726
rect 66100 19390 66186 19442
rect 66238 19390 66324 19442
rect 66100 19106 66324 19390
rect 66100 19054 66186 19106
rect 66238 19054 66324 19106
rect 66100 18772 66324 19054
rect 66100 18716 66184 18772
rect 66240 18716 66324 18772
rect 66100 18434 66324 18716
rect 66100 18382 66186 18434
rect 66238 18382 66324 18434
rect 66100 18098 66324 18382
rect 66100 18046 66186 18098
rect 66238 18046 66324 18098
rect 66100 17762 66324 18046
rect 66100 17710 66186 17762
rect 66238 17710 66324 17762
rect 66100 17426 66324 17710
rect 66100 17374 66186 17426
rect 66238 17374 66324 17426
rect 66100 17092 66324 17374
rect 66100 17036 66184 17092
rect 66240 17036 66324 17092
rect 66100 16754 66324 17036
rect 66100 16702 66186 16754
rect 66238 16702 66324 16754
rect 66100 16418 66324 16702
rect 66100 16366 66186 16418
rect 66238 16366 66324 16418
rect 66100 16082 66324 16366
rect 66100 16030 66186 16082
rect 66238 16030 66324 16082
rect 66100 15746 66324 16030
rect 66100 15694 66186 15746
rect 66238 15694 66324 15746
rect 66100 15412 66324 15694
rect 66100 15356 66184 15412
rect 66240 15356 66324 15412
rect 66100 15074 66324 15356
rect 66100 15022 66186 15074
rect 66238 15022 66324 15074
rect 66100 14738 66324 15022
rect 66100 14686 66186 14738
rect 66238 14686 66324 14738
rect 66100 14402 66324 14686
rect 56872 14368 56928 14377
rect 18442 13014 18470 14349
rect 56872 14303 56928 14312
rect 66100 14350 66186 14402
rect 66238 14350 66324 14402
rect 57954 14112 58010 14121
rect 56671 14041 56727 14050
rect 56671 13976 56727 13985
rect 57009 14041 57065 14050
rect 57954 14047 58010 14056
rect 66100 14066 66324 14350
rect 57009 13976 57065 13985
rect 66100 14014 66186 14066
rect 66238 14014 66324 14066
rect 18428 13005 18484 13014
rect 18428 12940 18484 12949
rect 21469 10186 21497 13822
rect 66100 13732 66324 14014
rect 66100 13676 66184 13732
rect 66240 13676 66324 13732
rect 66100 13394 66324 13676
rect 66100 13342 66186 13394
rect 66238 13342 66324 13394
rect 66100 13058 66324 13342
rect 66100 13006 66186 13058
rect 66238 13006 66324 13058
rect 66100 12722 66324 13006
rect 66100 12670 66186 12722
rect 66238 12670 66324 12722
rect 56591 12483 56647 12492
rect 56591 12418 56647 12427
rect 57009 12483 57065 12492
rect 57009 12418 57065 12427
rect 57954 12412 58010 12421
rect 57954 12347 58010 12356
rect 66100 12386 66324 12670
rect 66100 12334 66186 12386
rect 66238 12334 66324 12386
rect 66100 12052 66324 12334
rect 66100 11996 66184 12052
rect 66240 11996 66324 12052
rect 66100 11714 66324 11996
rect 66100 11662 66186 11714
rect 66238 11662 66324 11714
rect 66100 11378 66324 11662
rect 66100 11326 66186 11378
rect 66238 11326 66324 11378
rect 57954 11284 58010 11293
rect 56511 11213 56567 11222
rect 56511 11148 56567 11157
rect 57009 11213 57065 11222
rect 57954 11219 58010 11228
rect 57009 11148 57065 11157
rect 66100 11042 66324 11326
rect 66100 10990 66186 11042
rect 66238 10990 66324 11042
rect 66100 10706 66324 10990
rect 66100 10654 66186 10706
rect 66238 10654 66324 10706
rect 66100 10372 66324 10654
rect 66100 10316 66184 10372
rect 66240 10316 66324 10372
rect 21455 10177 21511 10186
rect 21455 10112 21511 10121
rect 66100 10034 66324 10316
rect 66100 9982 66186 10034
rect 66238 9982 66324 10034
rect 66100 9698 66324 9982
rect 56431 9655 56487 9664
rect 56431 9590 56487 9599
rect 57009 9655 57065 9664
rect 57009 9590 57065 9599
rect 66100 9646 66186 9698
rect 66238 9646 66324 9698
rect 57954 9584 58010 9593
rect 57954 9519 58010 9528
rect 66100 9362 66324 9646
rect 66100 9310 66186 9362
rect 66238 9310 66324 9362
rect 66100 9026 66324 9310
rect 66100 8974 66186 9026
rect 66238 8974 66324 9026
rect 21579 8763 21635 8772
rect 21579 8698 21635 8707
rect 21593 6370 21621 8698
rect 66100 8692 66324 8974
rect 66100 8636 66184 8692
rect 66240 8636 66324 8692
rect 57954 8456 58010 8465
rect 56351 8385 56407 8394
rect 56351 8320 56407 8329
rect 57009 8385 57065 8394
rect 57954 8391 58010 8400
rect 57009 8320 57065 8329
rect 66100 8354 66324 8636
rect 66100 8302 66186 8354
rect 66238 8302 66324 8354
rect 66100 8018 66324 8302
rect 66100 7966 66186 8018
rect 66238 7966 66324 8018
rect 66100 7682 66324 7966
rect 66100 7630 66186 7682
rect 66238 7630 66324 7682
rect 66100 7346 66324 7630
rect 66100 7294 66186 7346
rect 66238 7294 66324 7346
rect 66100 7012 66324 7294
rect 66100 6956 66184 7012
rect 66240 6956 66324 7012
rect 56271 6827 56327 6836
rect 56271 6762 56327 6771
rect 57009 6827 57065 6836
rect 57009 6762 57065 6771
rect 57954 6756 58010 6765
rect 57954 6691 58010 6700
rect 66100 6674 66324 6956
rect 66100 6622 66186 6674
rect 66238 6622 66324 6674
rect 6005 4483 6061 4492
rect 10836 4479 10934 4507
rect 6005 4418 6061 4427
rect 1496 4270 1582 4322
rect 1634 4270 1720 4322
rect 2708 4378 2764 4387
rect 2708 4313 2764 4322
rect 1496 3986 1720 4270
rect 1496 3934 1582 3986
rect 1634 3934 1720 3986
rect 1496 3652 1720 3934
rect 1496 3596 1580 3652
rect 1636 3596 1720 3652
rect 1496 3314 1720 3596
rect 1496 3262 1582 3314
rect 1634 3262 1720 3314
rect 1496 2978 1720 3262
rect 1496 2926 1582 2978
rect 1634 2926 1720 2978
rect 1496 2642 1720 2926
rect 10906 2793 10934 4479
rect 66100 6338 66324 6622
rect 66100 6286 66186 6338
rect 66238 6286 66324 6338
rect 66100 6002 66324 6286
rect 66100 5950 66186 6002
rect 66238 5950 66324 6002
rect 66100 5666 66324 5950
rect 66100 5614 66186 5666
rect 66238 5614 66324 5666
rect 66100 5332 66324 5614
rect 66100 5276 66184 5332
rect 66240 5276 66324 5332
rect 66100 4994 66324 5276
rect 66100 4942 66186 4994
rect 66238 4942 66324 4994
rect 66100 4658 66324 4942
rect 66100 4606 66186 4658
rect 66238 4606 66324 4658
rect 66100 4322 66324 4606
rect 66100 4270 66186 4322
rect 66238 4270 66324 4322
rect 66100 3986 66324 4270
rect 66100 3934 66186 3986
rect 66238 3934 66324 3986
rect 66100 3652 66324 3934
rect 66100 3596 66184 3652
rect 66240 3596 66324 3652
rect 66100 3314 66324 3596
rect 66100 3262 66186 3314
rect 66238 3262 66324 3314
rect 12146 3040 12202 3049
rect 12146 2975 12202 2984
rect 13314 3040 13370 3049
rect 13314 2975 13370 2984
rect 14482 3040 14538 3049
rect 14482 2975 14538 2984
rect 15650 3040 15706 3049
rect 15650 2975 15706 2984
rect 16818 3040 16874 3049
rect 16818 2975 16874 2984
rect 17986 3040 18042 3049
rect 17986 2975 18042 2984
rect 19154 3040 19210 3049
rect 19154 2975 19210 2984
rect 20322 3040 20378 3049
rect 20322 2975 20378 2984
rect 21490 3040 21546 3049
rect 21490 2975 21546 2984
rect 22658 3040 22714 3049
rect 22658 2975 22714 2984
rect 66100 2978 66324 3262
rect 66100 2926 66186 2978
rect 66238 2926 66324 2978
rect 10892 2784 10948 2793
rect 10892 2719 10948 2728
rect 1496 2590 1582 2642
rect 1634 2590 1720 2642
rect 1496 2306 1720 2590
rect 1496 2254 1582 2306
rect 1634 2254 1720 2306
rect 1496 1972 1720 2254
rect 1496 1916 1580 1972
rect 1636 1916 1720 1972
rect 1496 1496 1720 1916
rect 66100 2642 66324 2926
rect 66100 2590 66186 2642
rect 66238 2590 66324 2642
rect 66100 2306 66324 2590
rect 66100 2254 66186 2306
rect 66238 2254 66324 2306
rect 66100 1972 66324 2254
rect 66100 1916 66184 1972
rect 66240 1916 66324 1972
rect 1916 1636 1972 1645
rect 1916 1571 1972 1580
rect 3596 1636 3652 1645
rect 3596 1571 3652 1580
rect 5276 1636 5332 1645
rect 5276 1571 5332 1580
rect 6956 1636 7012 1645
rect 6956 1571 7012 1580
rect 8636 1636 8692 1645
rect 8636 1571 8692 1580
rect 10316 1636 10372 1645
rect 10316 1571 10372 1580
rect 11996 1636 12052 1645
rect 11996 1571 12052 1580
rect 13676 1636 13732 1645
rect 13676 1571 13732 1580
rect 15356 1636 15412 1645
rect 15356 1571 15412 1580
rect 17036 1636 17092 1645
rect 17036 1571 17092 1580
rect 18716 1636 18772 1645
rect 18716 1571 18772 1580
rect 20396 1636 20452 1645
rect 20396 1571 20452 1580
rect 22076 1636 22132 1645
rect 22076 1571 22132 1580
rect 23756 1636 23812 1645
rect 23756 1571 23812 1580
rect 25436 1636 25492 1645
rect 25436 1571 25492 1580
rect 27116 1636 27172 1645
rect 27116 1571 27172 1580
rect 28796 1636 28852 1645
rect 28796 1571 28852 1580
rect 30476 1636 30532 1645
rect 30476 1571 30532 1580
rect 32156 1636 32212 1645
rect 32156 1571 32212 1580
rect 33836 1636 33892 1645
rect 33836 1571 33892 1580
rect 35516 1636 35572 1645
rect 35516 1571 35572 1580
rect 37196 1636 37252 1645
rect 37196 1571 37252 1580
rect 38876 1636 38932 1645
rect 38876 1571 38932 1580
rect 40556 1636 40612 1645
rect 40556 1571 40612 1580
rect 42236 1636 42292 1645
rect 42236 1571 42292 1580
rect 43916 1636 43972 1645
rect 43916 1571 43972 1580
rect 45596 1636 45652 1645
rect 45596 1571 45652 1580
rect 47276 1636 47332 1645
rect 47276 1571 47332 1580
rect 48956 1636 49012 1645
rect 48956 1571 49012 1580
rect 50636 1636 50692 1645
rect 50636 1571 50692 1580
rect 52316 1636 52372 1645
rect 52316 1571 52372 1580
rect 53996 1636 54052 1645
rect 53996 1571 54052 1580
rect 55676 1636 55732 1645
rect 55676 1571 55732 1580
rect 57356 1636 57412 1645
rect 57356 1571 57412 1580
rect 59036 1636 59092 1645
rect 59036 1571 59092 1580
rect 60716 1636 60772 1645
rect 60716 1571 60772 1580
rect 62396 1636 62452 1645
rect 62396 1571 62452 1580
rect 64076 1636 64132 1645
rect 64076 1571 64132 1580
rect 65756 1636 65812 1645
rect 65756 1571 65812 1580
rect 66100 1496 66324 1916
<< via2 >>
rect 1916 51156 1972 51158
rect 1916 51104 1918 51156
rect 1918 51104 1970 51156
rect 1970 51104 1972 51156
rect 1916 51102 1972 51104
rect 3596 51156 3652 51158
rect 3596 51104 3598 51156
rect 3598 51104 3650 51156
rect 3650 51104 3652 51156
rect 3596 51102 3652 51104
rect 5276 51156 5332 51158
rect 5276 51104 5278 51156
rect 5278 51104 5330 51156
rect 5330 51104 5332 51156
rect 5276 51102 5332 51104
rect 6956 51156 7012 51158
rect 6956 51104 6958 51156
rect 6958 51104 7010 51156
rect 7010 51104 7012 51156
rect 6956 51102 7012 51104
rect 8636 51156 8692 51158
rect 8636 51104 8638 51156
rect 8638 51104 8690 51156
rect 8690 51104 8692 51156
rect 8636 51102 8692 51104
rect 10316 51156 10372 51158
rect 10316 51104 10318 51156
rect 10318 51104 10370 51156
rect 10370 51104 10372 51156
rect 10316 51102 10372 51104
rect 11996 51156 12052 51158
rect 11996 51104 11998 51156
rect 11998 51104 12050 51156
rect 12050 51104 12052 51156
rect 11996 51102 12052 51104
rect 13676 51156 13732 51158
rect 13676 51104 13678 51156
rect 13678 51104 13730 51156
rect 13730 51104 13732 51156
rect 13676 51102 13732 51104
rect 15356 51156 15412 51158
rect 15356 51104 15358 51156
rect 15358 51104 15410 51156
rect 15410 51104 15412 51156
rect 15356 51102 15412 51104
rect 17036 51156 17092 51158
rect 17036 51104 17038 51156
rect 17038 51104 17090 51156
rect 17090 51104 17092 51156
rect 17036 51102 17092 51104
rect 18716 51156 18772 51158
rect 18716 51104 18718 51156
rect 18718 51104 18770 51156
rect 18770 51104 18772 51156
rect 18716 51102 18772 51104
rect 20396 51156 20452 51158
rect 20396 51104 20398 51156
rect 20398 51104 20450 51156
rect 20450 51104 20452 51156
rect 20396 51102 20452 51104
rect 22076 51156 22132 51158
rect 22076 51104 22078 51156
rect 22078 51104 22130 51156
rect 22130 51104 22132 51156
rect 22076 51102 22132 51104
rect 23756 51156 23812 51158
rect 23756 51104 23758 51156
rect 23758 51104 23810 51156
rect 23810 51104 23812 51156
rect 23756 51102 23812 51104
rect 25436 51156 25492 51158
rect 25436 51104 25438 51156
rect 25438 51104 25490 51156
rect 25490 51104 25492 51156
rect 25436 51102 25492 51104
rect 27116 51156 27172 51158
rect 27116 51104 27118 51156
rect 27118 51104 27170 51156
rect 27170 51104 27172 51156
rect 27116 51102 27172 51104
rect 28796 51156 28852 51158
rect 28796 51104 28798 51156
rect 28798 51104 28850 51156
rect 28850 51104 28852 51156
rect 28796 51102 28852 51104
rect 30476 51156 30532 51158
rect 30476 51104 30478 51156
rect 30478 51104 30530 51156
rect 30530 51104 30532 51156
rect 30476 51102 30532 51104
rect 32156 51156 32212 51158
rect 32156 51104 32158 51156
rect 32158 51104 32210 51156
rect 32210 51104 32212 51156
rect 32156 51102 32212 51104
rect 33836 51156 33892 51158
rect 33836 51104 33838 51156
rect 33838 51104 33890 51156
rect 33890 51104 33892 51156
rect 33836 51102 33892 51104
rect 35516 51156 35572 51158
rect 35516 51104 35518 51156
rect 35518 51104 35570 51156
rect 35570 51104 35572 51156
rect 35516 51102 35572 51104
rect 37196 51156 37252 51158
rect 37196 51104 37198 51156
rect 37198 51104 37250 51156
rect 37250 51104 37252 51156
rect 37196 51102 37252 51104
rect 38876 51156 38932 51158
rect 38876 51104 38878 51156
rect 38878 51104 38930 51156
rect 38930 51104 38932 51156
rect 38876 51102 38932 51104
rect 40556 51156 40612 51158
rect 40556 51104 40558 51156
rect 40558 51104 40610 51156
rect 40610 51104 40612 51156
rect 40556 51102 40612 51104
rect 42236 51156 42292 51158
rect 42236 51104 42238 51156
rect 42238 51104 42290 51156
rect 42290 51104 42292 51156
rect 42236 51102 42292 51104
rect 43916 51156 43972 51158
rect 43916 51104 43918 51156
rect 43918 51104 43970 51156
rect 43970 51104 43972 51156
rect 43916 51102 43972 51104
rect 45596 51156 45652 51158
rect 45596 51104 45598 51156
rect 45598 51104 45650 51156
rect 45650 51104 45652 51156
rect 45596 51102 45652 51104
rect 47276 51156 47332 51158
rect 47276 51104 47278 51156
rect 47278 51104 47330 51156
rect 47330 51104 47332 51156
rect 47276 51102 47332 51104
rect 48956 51156 49012 51158
rect 48956 51104 48958 51156
rect 48958 51104 49010 51156
rect 49010 51104 49012 51156
rect 48956 51102 49012 51104
rect 50636 51156 50692 51158
rect 50636 51104 50638 51156
rect 50638 51104 50690 51156
rect 50690 51104 50692 51156
rect 50636 51102 50692 51104
rect 52316 51156 52372 51158
rect 52316 51104 52318 51156
rect 52318 51104 52370 51156
rect 52370 51104 52372 51156
rect 52316 51102 52372 51104
rect 53996 51156 54052 51158
rect 53996 51104 53998 51156
rect 53998 51104 54050 51156
rect 54050 51104 54052 51156
rect 53996 51102 54052 51104
rect 55676 51156 55732 51158
rect 55676 51104 55678 51156
rect 55678 51104 55730 51156
rect 55730 51104 55732 51156
rect 55676 51102 55732 51104
rect 57356 51156 57412 51158
rect 57356 51104 57358 51156
rect 57358 51104 57410 51156
rect 57410 51104 57412 51156
rect 57356 51102 57412 51104
rect 59036 51156 59092 51158
rect 59036 51104 59038 51156
rect 59038 51104 59090 51156
rect 59090 51104 59092 51156
rect 59036 51102 59092 51104
rect 60716 51156 60772 51158
rect 60716 51104 60718 51156
rect 60718 51104 60770 51156
rect 60770 51104 60772 51156
rect 60716 51102 60772 51104
rect 62396 51156 62452 51158
rect 62396 51104 62398 51156
rect 62398 51104 62450 51156
rect 62450 51104 62452 51156
rect 62396 51102 62452 51104
rect 64076 51156 64132 51158
rect 64076 51104 64078 51156
rect 64078 51104 64130 51156
rect 64130 51104 64132 51156
rect 64076 51102 64132 51104
rect 65756 51156 65812 51158
rect 65756 51104 65758 51156
rect 65758 51104 65810 51156
rect 65810 51104 65812 51156
rect 65756 51102 65812 51104
rect 1580 50690 1636 50692
rect 1580 50638 1582 50690
rect 1582 50638 1634 50690
rect 1634 50638 1636 50690
rect 1580 50636 1636 50638
rect 66184 50690 66240 50692
rect 66184 50638 66186 50690
rect 66186 50638 66238 50690
rect 66238 50638 66240 50690
rect 66184 50636 66240 50638
rect 56872 49954 56928 50010
rect 53282 49698 53338 49754
rect 54450 49698 54506 49754
rect 1580 49010 1636 49012
rect 1580 48958 1582 49010
rect 1582 48958 1634 49010
rect 1634 48958 1636 49010
rect 1580 48956 1636 48958
rect 1580 47330 1636 47332
rect 1580 47278 1582 47330
rect 1582 47278 1634 47330
rect 1634 47278 1636 47330
rect 1580 47276 1636 47278
rect 66184 49010 66240 49012
rect 66184 48958 66186 49010
rect 66186 48958 66238 49010
rect 66238 48958 66240 49010
rect 66184 48956 66240 48958
rect 65056 48734 65112 48790
rect 61759 48629 61815 48685
rect 23983 46887 24039 46889
rect 23983 46835 23985 46887
rect 23985 46835 24037 46887
rect 24037 46835 24039 46887
rect 23983 46833 24039 46835
rect 26479 46887 26535 46889
rect 26479 46835 26481 46887
rect 26481 46835 26533 46887
rect 26533 46835 26535 46887
rect 26479 46833 26535 46835
rect 28975 46887 29031 46889
rect 28975 46835 28977 46887
rect 28977 46835 29029 46887
rect 29029 46835 29031 46887
rect 28975 46833 29031 46835
rect 31471 46887 31527 46889
rect 31471 46835 31473 46887
rect 31473 46835 31525 46887
rect 31525 46835 31527 46887
rect 31471 46833 31527 46835
rect 33967 46887 34023 46889
rect 33967 46835 33969 46887
rect 33969 46835 34021 46887
rect 34021 46835 34023 46887
rect 33967 46833 34023 46835
rect 36463 46887 36519 46889
rect 36463 46835 36465 46887
rect 36465 46835 36517 46887
rect 36517 46835 36519 46887
rect 36463 46833 36519 46835
rect 38959 46887 39015 46889
rect 38959 46835 38961 46887
rect 38961 46835 39013 46887
rect 39013 46835 39015 46887
rect 38959 46833 39015 46835
rect 41455 46887 41511 46889
rect 41455 46835 41457 46887
rect 41457 46835 41509 46887
rect 41509 46835 41511 46887
rect 41455 46833 41511 46835
rect 1580 45650 1636 45652
rect 1580 45598 1582 45650
rect 1582 45598 1634 45650
rect 1634 45598 1636 45650
rect 1580 45596 1636 45598
rect 46067 44333 46123 44389
rect 1580 43970 1636 43972
rect 1580 43918 1582 43970
rect 1582 43918 1634 43970
rect 1634 43918 1636 43970
rect 1580 43916 1636 43918
rect 1580 42290 1636 42292
rect 1580 42238 1582 42290
rect 1582 42238 1634 42290
rect 1634 42238 1636 42290
rect 1580 42236 1636 42238
rect 46191 42935 46247 42991
rect 49252 41521 49308 41577
rect 1580 40610 1636 40612
rect 1580 40558 1582 40610
rect 1582 40558 1634 40610
rect 1634 40558 1636 40610
rect 1580 40556 1636 40558
rect 46769 40152 46825 40153
rect 46769 40100 46771 40152
rect 46771 40100 46823 40152
rect 46823 40100 46825 40152
rect 46769 40097 46825 40100
rect 48660 40139 48716 40141
rect 48660 40087 48662 40139
rect 48662 40087 48714 40139
rect 48714 40087 48716 40139
rect 48660 40085 48716 40087
rect 1580 38930 1636 38932
rect 1580 38878 1582 38930
rect 1582 38878 1634 38930
rect 1634 38878 1636 38930
rect 1580 38876 1636 38878
rect 1580 37250 1636 37252
rect 1580 37198 1582 37250
rect 1582 37198 1634 37250
rect 1634 37198 1636 37250
rect 1580 37196 1636 37198
rect 1580 35570 1636 35572
rect 1580 35518 1582 35570
rect 1582 35518 1634 35570
rect 1634 35518 1636 35570
rect 1580 35516 1636 35518
rect 1580 33890 1636 33892
rect 1580 33838 1582 33890
rect 1582 33838 1634 33890
rect 1634 33838 1636 33890
rect 1580 33836 1636 33838
rect 1580 32210 1636 32212
rect 1580 32158 1582 32210
rect 1582 32158 1634 32210
rect 1634 32158 1636 32210
rect 1580 32156 1636 32158
rect 1580 30530 1636 30532
rect 1580 30478 1582 30530
rect 1582 30478 1634 30530
rect 1634 30478 1636 30530
rect 1580 30476 1636 30478
rect 9810 30220 9866 30276
rect 10755 30149 10811 30205
rect 11409 30203 11465 30205
rect 11409 30151 11411 30203
rect 11411 30151 11463 30203
rect 11463 30151 11465 30203
rect 11409 30149 11465 30151
rect 1580 28850 1636 28852
rect 1580 28798 1582 28850
rect 1582 28798 1634 28850
rect 1634 28798 1636 28850
rect 1580 28796 1636 28798
rect 10755 28591 10811 28647
rect 11329 28645 11385 28647
rect 11329 28593 11331 28645
rect 11331 28593 11383 28645
rect 11383 28593 11385 28645
rect 11329 28591 11385 28593
rect 9810 28520 9866 28576
rect 9810 27392 9866 27448
rect 10755 27321 10811 27377
rect 11249 27375 11305 27377
rect 11249 27323 11251 27375
rect 11251 27323 11303 27375
rect 11303 27323 11305 27375
rect 11249 27321 11305 27323
rect 1580 27170 1636 27172
rect 1580 27118 1582 27170
rect 1582 27118 1634 27170
rect 1634 27118 1636 27170
rect 1580 27116 1636 27118
rect 10755 25763 10811 25819
rect 11169 25817 11225 25819
rect 11169 25765 11171 25817
rect 11171 25765 11223 25817
rect 11223 25765 11225 25817
rect 11169 25763 11225 25765
rect 9810 25692 9866 25748
rect 1580 25490 1636 25492
rect 1580 25438 1582 25490
rect 1582 25438 1634 25490
rect 1634 25438 1636 25490
rect 1580 25436 1636 25438
rect 9810 24564 9866 24620
rect 10755 24493 10811 24549
rect 11089 24547 11145 24549
rect 11089 24495 11091 24547
rect 11091 24495 11143 24547
rect 11143 24495 11145 24547
rect 11089 24493 11145 24495
rect 1580 23810 1636 23812
rect 1580 23758 1582 23810
rect 1582 23758 1634 23810
rect 1634 23758 1636 23810
rect 1580 23756 1636 23758
rect 10755 22935 10811 22991
rect 11009 22989 11065 22991
rect 11009 22937 11011 22989
rect 11011 22937 11063 22989
rect 11063 22937 11065 22989
rect 11009 22935 11065 22937
rect 9810 22864 9866 22920
rect 10892 22608 10948 22664
rect 1580 22130 1636 22132
rect 1580 22078 1582 22130
rect 1582 22078 1634 22130
rect 1634 22078 1636 22130
rect 1580 22076 1636 22078
rect 2495 21471 2551 21527
rect 1580 20450 1636 20452
rect 1580 20398 1582 20450
rect 1582 20398 1634 20450
rect 1634 20398 1636 20450
rect 1580 20396 1636 20398
rect 1580 18770 1636 18772
rect 1580 18718 1582 18770
rect 1582 18718 1634 18770
rect 1634 18718 1636 18770
rect 1580 18716 1636 18718
rect 1580 17090 1636 17092
rect 1580 17038 1582 17090
rect 1582 17038 1634 17090
rect 1634 17038 1636 17090
rect 1580 17036 1636 17038
rect 1580 15410 1636 15412
rect 1580 15358 1582 15410
rect 1582 15358 1634 15410
rect 1634 15358 1636 15410
rect 1580 15356 1636 15358
rect 1580 13730 1636 13732
rect 1580 13678 1582 13730
rect 1582 13678 1634 13730
rect 1634 13678 1636 13730
rect 1580 13676 1636 13678
rect 10808 12949 10864 13005
rect 1580 12050 1636 12052
rect 1580 11998 1582 12050
rect 1582 11998 1634 12050
rect 1634 11998 1636 12050
rect 1580 11996 1636 11998
rect 1580 10370 1636 10372
rect 1580 10318 1582 10370
rect 1582 10318 1634 10370
rect 1634 10318 1636 10370
rect 1580 10316 1636 10318
rect 10808 10121 10864 10177
rect 10808 8707 10864 8763
rect 1580 8690 1636 8692
rect 1580 8638 1582 8690
rect 1582 8638 1634 8690
rect 1634 8638 1636 8690
rect 1580 8636 1636 8638
rect 1580 7010 1636 7012
rect 1580 6958 1582 7010
rect 1582 6958 1634 7010
rect 1634 6958 1636 7010
rect 1580 6956 1636 6958
rect 1580 5330 1636 5332
rect 1580 5278 1582 5330
rect 1582 5278 1634 5330
rect 1634 5278 1636 5330
rect 1580 5276 1636 5278
rect 19020 14489 19076 14491
rect 19020 14437 19022 14489
rect 19022 14437 19074 14489
rect 19074 14437 19076 14489
rect 19020 14435 19076 14437
rect 20911 14476 20967 14479
rect 20911 14424 20913 14476
rect 20913 14424 20965 14476
rect 20965 14424 20967 14476
rect 20911 14423 20967 14424
rect 66184 47330 66240 47332
rect 66184 47278 66186 47330
rect 66186 47278 66238 47330
rect 66238 47278 66240 47330
rect 66184 47276 66240 47278
rect 66184 45650 66240 45652
rect 66184 45598 66186 45650
rect 66186 45598 66238 45650
rect 66238 45598 66240 45650
rect 66184 45596 66240 45598
rect 56956 44333 57012 44389
rect 66184 43970 66240 43972
rect 66184 43918 66186 43970
rect 66186 43918 66238 43970
rect 66238 43918 66240 43970
rect 66184 43916 66240 43918
rect 56956 42935 57012 42991
rect 66184 42290 66240 42292
rect 66184 42238 66186 42290
rect 66186 42238 66238 42290
rect 66238 42238 66240 42290
rect 66184 42236 66240 42238
rect 56956 41521 57012 41577
rect 66184 40610 66240 40612
rect 66184 40558 66186 40610
rect 66186 40558 66238 40610
rect 66238 40558 66240 40610
rect 66184 40556 66240 40558
rect 66184 38930 66240 38932
rect 66184 38878 66186 38930
rect 66186 38878 66238 38930
rect 66238 38878 66240 38930
rect 66184 38876 66240 38878
rect 66184 37250 66240 37252
rect 66184 37198 66186 37250
rect 66186 37198 66238 37250
rect 66238 37198 66240 37250
rect 66184 37196 66240 37198
rect 66184 35570 66240 35572
rect 66184 35518 66186 35570
rect 66186 35518 66238 35570
rect 66238 35518 66240 35570
rect 66184 35516 66240 35518
rect 66184 33890 66240 33892
rect 66184 33838 66186 33890
rect 66186 33838 66238 33890
rect 66238 33838 66240 33890
rect 66184 33836 66240 33838
rect 66184 32210 66240 32212
rect 66184 32158 66186 32210
rect 66186 32158 66238 32210
rect 66238 32158 66240 32210
rect 66184 32156 66240 32158
rect 65269 31585 65325 31641
rect 66184 30530 66240 30532
rect 66184 30478 66186 30530
rect 66186 30478 66238 30530
rect 66238 30478 66240 30530
rect 66184 30476 66240 30478
rect 66184 28850 66240 28852
rect 66184 28798 66186 28850
rect 66186 28798 66238 28850
rect 66238 28798 66240 28850
rect 66184 28796 66240 28798
rect 66184 27170 66240 27172
rect 66184 27118 66186 27170
rect 66186 27118 66238 27170
rect 66238 27118 66240 27170
rect 66184 27116 66240 27118
rect 66184 25490 66240 25492
rect 66184 25438 66186 25490
rect 66186 25438 66238 25490
rect 66238 25438 66240 25490
rect 66184 25436 66240 25438
rect 66184 23810 66240 23812
rect 66184 23758 66186 23810
rect 66186 23758 66238 23810
rect 66238 23758 66240 23810
rect 66184 23756 66240 23758
rect 66184 22130 66240 22132
rect 66184 22078 66186 22130
rect 66186 22078 66238 22130
rect 66238 22078 66240 22130
rect 66184 22076 66240 22078
rect 66184 20450 66240 20452
rect 66184 20398 66186 20450
rect 66186 20398 66238 20450
rect 66238 20398 66240 20450
rect 66184 20396 66240 20398
rect 66184 18770 66240 18772
rect 66184 18718 66186 18770
rect 66186 18718 66238 18770
rect 66238 18718 66240 18770
rect 66184 18716 66240 18718
rect 66184 17090 66240 17092
rect 66184 17038 66186 17090
rect 66186 17038 66238 17090
rect 66238 17038 66240 17090
rect 66184 17036 66240 17038
rect 66184 15410 66240 15412
rect 66184 15358 66186 15410
rect 66186 15358 66238 15410
rect 66238 15358 66240 15410
rect 66184 15356 66240 15358
rect 56872 14312 56928 14368
rect 57954 14056 58010 14112
rect 56671 14039 56727 14041
rect 56671 13987 56673 14039
rect 56673 13987 56725 14039
rect 56725 13987 56727 14039
rect 56671 13985 56727 13987
rect 57009 13985 57065 14041
rect 18428 12949 18484 13005
rect 66184 13730 66240 13732
rect 66184 13678 66186 13730
rect 66186 13678 66238 13730
rect 66238 13678 66240 13730
rect 66184 13676 66240 13678
rect 56591 12481 56647 12483
rect 56591 12429 56593 12481
rect 56593 12429 56645 12481
rect 56645 12429 56647 12481
rect 56591 12427 56647 12429
rect 57009 12427 57065 12483
rect 57954 12356 58010 12412
rect 66184 12050 66240 12052
rect 66184 11998 66186 12050
rect 66186 11998 66238 12050
rect 66238 11998 66240 12050
rect 66184 11996 66240 11998
rect 57954 11228 58010 11284
rect 56511 11211 56567 11213
rect 56511 11159 56513 11211
rect 56513 11159 56565 11211
rect 56565 11159 56567 11211
rect 56511 11157 56567 11159
rect 57009 11157 57065 11213
rect 66184 10370 66240 10372
rect 66184 10318 66186 10370
rect 66186 10318 66238 10370
rect 66238 10318 66240 10370
rect 66184 10316 66240 10318
rect 21455 10121 21511 10177
rect 56431 9653 56487 9655
rect 56431 9601 56433 9653
rect 56433 9601 56485 9653
rect 56485 9601 56487 9653
rect 56431 9599 56487 9601
rect 57009 9599 57065 9655
rect 57954 9528 58010 9584
rect 21579 8707 21635 8763
rect 66184 8690 66240 8692
rect 66184 8638 66186 8690
rect 66186 8638 66238 8690
rect 66238 8638 66240 8690
rect 66184 8636 66240 8638
rect 57954 8400 58010 8456
rect 56351 8383 56407 8385
rect 56351 8331 56353 8383
rect 56353 8331 56405 8383
rect 56405 8331 56407 8383
rect 56351 8329 56407 8331
rect 57009 8329 57065 8385
rect 66184 7010 66240 7012
rect 66184 6958 66186 7010
rect 66186 6958 66238 7010
rect 66238 6958 66240 7010
rect 66184 6956 66240 6958
rect 56271 6825 56327 6827
rect 56271 6773 56273 6825
rect 56273 6773 56325 6825
rect 56325 6773 56327 6825
rect 56271 6771 56327 6773
rect 57009 6771 57065 6827
rect 57954 6700 58010 6756
rect 6005 4427 6061 4483
rect 2708 4322 2764 4378
rect 1580 3650 1636 3652
rect 1580 3598 1582 3650
rect 1582 3598 1634 3650
rect 1634 3598 1636 3650
rect 1580 3596 1636 3598
rect 66184 5330 66240 5332
rect 66184 5278 66186 5330
rect 66186 5278 66238 5330
rect 66238 5278 66240 5330
rect 66184 5276 66240 5278
rect 66184 3650 66240 3652
rect 66184 3598 66186 3650
rect 66186 3598 66238 3650
rect 66238 3598 66240 3650
rect 66184 3596 66240 3598
rect 12146 2984 12202 3040
rect 13314 2984 13370 3040
rect 14482 2984 14538 3040
rect 15650 2984 15706 3040
rect 16818 2984 16874 3040
rect 17986 2984 18042 3040
rect 19154 2984 19210 3040
rect 20322 2984 20378 3040
rect 21490 2984 21546 3040
rect 22658 2984 22714 3040
rect 10892 2728 10948 2784
rect 1580 1970 1636 1972
rect 1580 1918 1582 1970
rect 1582 1918 1634 1970
rect 1634 1918 1636 1970
rect 1580 1916 1636 1918
rect 66184 1970 66240 1972
rect 66184 1918 66186 1970
rect 66186 1918 66238 1970
rect 66238 1918 66240 1970
rect 66184 1916 66240 1918
rect 1916 1634 1972 1636
rect 1916 1582 1918 1634
rect 1918 1582 1970 1634
rect 1970 1582 1972 1634
rect 1916 1580 1972 1582
rect 3596 1634 3652 1636
rect 3596 1582 3598 1634
rect 3598 1582 3650 1634
rect 3650 1582 3652 1634
rect 3596 1580 3652 1582
rect 5276 1634 5332 1636
rect 5276 1582 5278 1634
rect 5278 1582 5330 1634
rect 5330 1582 5332 1634
rect 5276 1580 5332 1582
rect 6956 1634 7012 1636
rect 6956 1582 6958 1634
rect 6958 1582 7010 1634
rect 7010 1582 7012 1634
rect 6956 1580 7012 1582
rect 8636 1634 8692 1636
rect 8636 1582 8638 1634
rect 8638 1582 8690 1634
rect 8690 1582 8692 1634
rect 8636 1580 8692 1582
rect 10316 1634 10372 1636
rect 10316 1582 10318 1634
rect 10318 1582 10370 1634
rect 10370 1582 10372 1634
rect 10316 1580 10372 1582
rect 11996 1634 12052 1636
rect 11996 1582 11998 1634
rect 11998 1582 12050 1634
rect 12050 1582 12052 1634
rect 11996 1580 12052 1582
rect 13676 1634 13732 1636
rect 13676 1582 13678 1634
rect 13678 1582 13730 1634
rect 13730 1582 13732 1634
rect 13676 1580 13732 1582
rect 15356 1634 15412 1636
rect 15356 1582 15358 1634
rect 15358 1582 15410 1634
rect 15410 1582 15412 1634
rect 15356 1580 15412 1582
rect 17036 1634 17092 1636
rect 17036 1582 17038 1634
rect 17038 1582 17090 1634
rect 17090 1582 17092 1634
rect 17036 1580 17092 1582
rect 18716 1634 18772 1636
rect 18716 1582 18718 1634
rect 18718 1582 18770 1634
rect 18770 1582 18772 1634
rect 18716 1580 18772 1582
rect 20396 1634 20452 1636
rect 20396 1582 20398 1634
rect 20398 1582 20450 1634
rect 20450 1582 20452 1634
rect 20396 1580 20452 1582
rect 22076 1634 22132 1636
rect 22076 1582 22078 1634
rect 22078 1582 22130 1634
rect 22130 1582 22132 1634
rect 22076 1580 22132 1582
rect 23756 1634 23812 1636
rect 23756 1582 23758 1634
rect 23758 1582 23810 1634
rect 23810 1582 23812 1634
rect 23756 1580 23812 1582
rect 25436 1634 25492 1636
rect 25436 1582 25438 1634
rect 25438 1582 25490 1634
rect 25490 1582 25492 1634
rect 25436 1580 25492 1582
rect 27116 1634 27172 1636
rect 27116 1582 27118 1634
rect 27118 1582 27170 1634
rect 27170 1582 27172 1634
rect 27116 1580 27172 1582
rect 28796 1634 28852 1636
rect 28796 1582 28798 1634
rect 28798 1582 28850 1634
rect 28850 1582 28852 1634
rect 28796 1580 28852 1582
rect 30476 1634 30532 1636
rect 30476 1582 30478 1634
rect 30478 1582 30530 1634
rect 30530 1582 30532 1634
rect 30476 1580 30532 1582
rect 32156 1634 32212 1636
rect 32156 1582 32158 1634
rect 32158 1582 32210 1634
rect 32210 1582 32212 1634
rect 32156 1580 32212 1582
rect 33836 1634 33892 1636
rect 33836 1582 33838 1634
rect 33838 1582 33890 1634
rect 33890 1582 33892 1634
rect 33836 1580 33892 1582
rect 35516 1634 35572 1636
rect 35516 1582 35518 1634
rect 35518 1582 35570 1634
rect 35570 1582 35572 1634
rect 35516 1580 35572 1582
rect 37196 1634 37252 1636
rect 37196 1582 37198 1634
rect 37198 1582 37250 1634
rect 37250 1582 37252 1634
rect 37196 1580 37252 1582
rect 38876 1634 38932 1636
rect 38876 1582 38878 1634
rect 38878 1582 38930 1634
rect 38930 1582 38932 1634
rect 38876 1580 38932 1582
rect 40556 1634 40612 1636
rect 40556 1582 40558 1634
rect 40558 1582 40610 1634
rect 40610 1582 40612 1634
rect 40556 1580 40612 1582
rect 42236 1634 42292 1636
rect 42236 1582 42238 1634
rect 42238 1582 42290 1634
rect 42290 1582 42292 1634
rect 42236 1580 42292 1582
rect 43916 1634 43972 1636
rect 43916 1582 43918 1634
rect 43918 1582 43970 1634
rect 43970 1582 43972 1634
rect 43916 1580 43972 1582
rect 45596 1634 45652 1636
rect 45596 1582 45598 1634
rect 45598 1582 45650 1634
rect 45650 1582 45652 1634
rect 45596 1580 45652 1582
rect 47276 1634 47332 1636
rect 47276 1582 47278 1634
rect 47278 1582 47330 1634
rect 47330 1582 47332 1634
rect 47276 1580 47332 1582
rect 48956 1634 49012 1636
rect 48956 1582 48958 1634
rect 48958 1582 49010 1634
rect 49010 1582 49012 1634
rect 48956 1580 49012 1582
rect 50636 1634 50692 1636
rect 50636 1582 50638 1634
rect 50638 1582 50690 1634
rect 50690 1582 50692 1634
rect 50636 1580 50692 1582
rect 52316 1634 52372 1636
rect 52316 1582 52318 1634
rect 52318 1582 52370 1634
rect 52370 1582 52372 1634
rect 52316 1580 52372 1582
rect 53996 1634 54052 1636
rect 53996 1582 53998 1634
rect 53998 1582 54050 1634
rect 54050 1582 54052 1634
rect 53996 1580 54052 1582
rect 55676 1634 55732 1636
rect 55676 1582 55678 1634
rect 55678 1582 55730 1634
rect 55730 1582 55732 1634
rect 55676 1580 55732 1582
rect 57356 1634 57412 1636
rect 57356 1582 57358 1634
rect 57358 1582 57410 1634
rect 57410 1582 57412 1634
rect 57356 1580 57412 1582
rect 59036 1634 59092 1636
rect 59036 1582 59038 1634
rect 59038 1582 59090 1634
rect 59090 1582 59092 1634
rect 59036 1580 59092 1582
rect 60716 1634 60772 1636
rect 60716 1582 60718 1634
rect 60718 1582 60770 1634
rect 60770 1582 60772 1634
rect 60716 1580 60772 1582
rect 62396 1634 62452 1636
rect 62396 1582 62398 1634
rect 62398 1582 62450 1634
rect 62450 1582 62452 1634
rect 62396 1580 62452 1582
rect 64076 1634 64132 1636
rect 64076 1582 64078 1634
rect 64078 1582 64130 1634
rect 64130 1582 64132 1634
rect 64076 1580 64132 1582
rect 65756 1634 65812 1636
rect 65756 1582 65758 1634
rect 65758 1582 65810 1634
rect 65810 1582 65812 1634
rect 65756 1580 65812 1582
<< metal3 >>
rect 0 52732 67820 52738
rect 0 52668 6 52732
rect 70 52668 142 52732
rect 206 52668 278 52732
rect 342 52668 67478 52732
rect 67542 52668 67614 52732
rect 67678 52668 67750 52732
rect 67814 52668 67820 52732
rect 0 52596 67820 52668
rect 0 52532 6 52596
rect 70 52532 142 52596
rect 206 52532 278 52596
rect 342 52532 67478 52596
rect 67542 52532 67614 52596
rect 67678 52532 67750 52596
rect 67814 52532 67820 52596
rect 0 52460 67820 52532
rect 0 52396 6 52460
rect 70 52396 142 52460
rect 206 52396 278 52460
rect 342 52396 13672 52460
rect 13736 52396 27112 52460
rect 27176 52396 40552 52460
rect 40616 52396 53992 52460
rect 54056 52396 67478 52460
rect 67542 52396 67614 52460
rect 67678 52396 67750 52460
rect 67814 52396 67820 52460
rect 0 52390 67820 52396
rect 696 52036 67124 52042
rect 696 51972 702 52036
rect 766 51972 838 52036
rect 902 51972 974 52036
rect 1038 51972 66782 52036
rect 66846 51972 66918 52036
rect 66982 51972 67054 52036
rect 67118 51972 67124 52036
rect 696 51900 67124 51972
rect 696 51836 702 51900
rect 766 51836 838 51900
rect 902 51836 974 51900
rect 1038 51836 66782 51900
rect 66846 51836 66918 51900
rect 66982 51836 67054 51900
rect 67118 51836 67124 51900
rect 696 51764 67124 51836
rect 696 51700 702 51764
rect 766 51700 838 51764
rect 902 51700 974 51764
rect 1038 51700 14136 51764
rect 14200 51700 27297 51764
rect 27361 51700 40414 51764
rect 40478 51700 53448 51764
rect 53512 51700 66782 51764
rect 66846 51700 66918 51764
rect 66982 51700 67054 51764
rect 67118 51700 67124 51764
rect 696 51694 67124 51700
rect 1895 51168 1993 51179
rect 3575 51168 3673 51179
rect 5255 51168 5353 51179
rect 6935 51168 7033 51179
rect 8615 51168 8713 51179
rect 10295 51168 10393 51179
rect 11975 51168 12073 51179
rect 13655 51168 13753 51179
rect 15335 51168 15433 51179
rect 17015 51168 17113 51179
rect 18695 51168 18793 51179
rect 20375 51168 20473 51179
rect 22055 51168 22153 51179
rect 23735 51168 23833 51179
rect 25415 51168 25513 51179
rect 27095 51168 27193 51179
rect 28775 51168 28873 51179
rect 30455 51168 30553 51179
rect 32135 51168 32233 51179
rect 33815 51168 33913 51179
rect 35495 51168 35593 51179
rect 37175 51168 37273 51179
rect 38855 51168 38953 51179
rect 40535 51168 40633 51179
rect 42215 51168 42313 51179
rect 43895 51168 43993 51179
rect 45575 51168 45673 51179
rect 47255 51168 47353 51179
rect 48935 51168 49033 51179
rect 50615 51168 50713 51179
rect 52295 51168 52393 51179
rect 53975 51168 54073 51179
rect 55655 51168 55753 51179
rect 57335 51168 57433 51179
rect 59015 51168 59113 51179
rect 60695 51168 60793 51179
rect 62375 51168 62473 51179
rect 64055 51168 64153 51179
rect 65735 51168 65833 51179
rect 1895 51162 66250 51168
rect 1895 51098 1912 51162
rect 1976 51158 13672 51162
rect 13736 51158 27112 51162
rect 27176 51158 40552 51162
rect 40616 51158 53992 51162
rect 1976 51102 3596 51158
rect 3652 51102 5276 51158
rect 5332 51102 6956 51158
rect 7012 51102 8636 51158
rect 8692 51102 10316 51158
rect 10372 51102 11996 51158
rect 12052 51102 13672 51158
rect 13736 51102 15356 51158
rect 15412 51102 17036 51158
rect 17092 51102 18716 51158
rect 18772 51102 20396 51158
rect 20452 51102 22076 51158
rect 22132 51102 23756 51158
rect 23812 51102 25436 51158
rect 25492 51102 27112 51158
rect 27176 51102 28796 51158
rect 28852 51102 30476 51158
rect 30532 51102 32156 51158
rect 32212 51102 33836 51158
rect 33892 51102 35516 51158
rect 35572 51102 37196 51158
rect 37252 51102 38876 51158
rect 38932 51102 40552 51158
rect 40616 51102 42236 51158
rect 42292 51102 43916 51158
rect 43972 51102 45596 51158
rect 45652 51102 47276 51158
rect 47332 51102 48956 51158
rect 49012 51102 50636 51158
rect 50692 51102 52316 51158
rect 52372 51102 53992 51158
rect 1976 51098 13672 51102
rect 13736 51098 27112 51102
rect 27176 51098 40552 51102
rect 40616 51098 53992 51102
rect 54056 51098 54616 51162
rect 54680 51158 66180 51162
rect 54680 51102 55676 51158
rect 55732 51102 57356 51158
rect 57412 51102 59036 51158
rect 59092 51102 60716 51158
rect 60772 51102 62396 51158
rect 62452 51102 64076 51158
rect 64132 51102 65756 51158
rect 65812 51102 66180 51158
rect 54680 51098 66180 51102
rect 66244 51098 66250 51162
rect 1895 51092 66250 51098
rect 1895 51081 1993 51092
rect 3575 51081 3673 51092
rect 5255 51081 5353 51092
rect 6935 51081 7033 51092
rect 8615 51081 8713 51092
rect 10295 51081 10393 51092
rect 11975 51081 12073 51092
rect 13655 51081 13753 51092
rect 15335 51081 15433 51092
rect 17015 51081 17113 51092
rect 18695 51081 18793 51092
rect 20375 51081 20473 51092
rect 22055 51081 22153 51092
rect 23735 51081 23833 51092
rect 25415 51081 25513 51092
rect 27095 51081 27193 51092
rect 28775 51081 28873 51092
rect 30455 51081 30553 51092
rect 32135 51081 32233 51092
rect 33815 51081 33913 51092
rect 35495 51081 35593 51092
rect 37175 51081 37273 51092
rect 38855 51081 38953 51092
rect 40535 51081 40633 51092
rect 42215 51081 42313 51092
rect 43895 51081 43993 51092
rect 45575 51081 45673 51092
rect 47255 51081 47353 51092
rect 48935 51081 49033 51092
rect 50615 51081 50713 51092
rect 52295 51081 52393 51092
rect 53975 51081 54073 51092
rect 55655 51081 55753 51092
rect 57335 51081 57433 51092
rect 59015 51081 59113 51092
rect 60695 51081 60793 51092
rect 62375 51081 62473 51092
rect 64055 51081 64153 51092
rect 65735 51081 65833 51092
rect 1559 50702 1657 50713
rect 1559 50696 1982 50702
rect 1559 50632 1576 50696
rect 1640 50632 1912 50696
rect 1976 50632 1982 50696
rect 1559 50626 1982 50632
rect 66163 50696 66261 50713
rect 66163 50632 66180 50696
rect 66244 50632 66261 50696
rect 1559 50615 1657 50626
rect 66163 50615 66261 50632
rect 53431 50328 53529 50339
rect 52220 50322 61906 50328
rect 52220 50258 52226 50322
rect 52290 50258 53448 50322
rect 53512 50258 61836 50322
rect 61900 50258 61906 50322
rect 52220 50252 61906 50258
rect 53431 50241 53529 50252
rect 56867 50012 56933 50015
rect 53480 50010 56933 50012
rect 53480 49954 56872 50010
rect 56928 49954 56933 50010
rect 53480 49952 56933 49954
rect 56867 49949 56933 49952
rect 53261 49758 53359 49775
rect 53261 49694 53278 49758
rect 53342 49694 53359 49758
rect 53261 49677 53359 49694
rect 54429 49758 54527 49775
rect 54429 49694 54446 49758
rect 54510 49694 54527 49758
rect 54429 49677 54527 49694
rect 63928 49364 64026 49375
rect 62011 49358 64026 49364
rect 62011 49294 62017 49358
rect 62081 49294 64026 49358
rect 62011 49288 64026 49294
rect 63928 49277 64026 49288
rect 1559 49016 1657 49033
rect 1559 48952 1576 49016
rect 1640 48952 1657 49016
rect 1559 48935 1657 48952
rect 66163 49016 66261 49033
rect 66163 48952 66180 49016
rect 66244 48952 66261 49016
rect 66163 48935 66261 48952
rect 54599 48914 54697 48925
rect 54599 48908 57106 48914
rect 54599 48844 54616 48908
rect 54680 48844 57036 48908
rect 57100 48844 57106 48908
rect 54599 48838 57106 48844
rect 61692 48838 61825 48844
rect 54599 48827 54697 48838
rect 61692 48774 61698 48838
rect 61762 48774 61825 48838
rect 61692 48768 61825 48774
rect 61749 48706 61825 48768
rect 65035 48800 65133 48811
rect 65035 48790 67820 48800
rect 65035 48734 65056 48790
rect 65112 48734 67820 48790
rect 65035 48724 67820 48734
rect 65035 48713 65133 48724
rect 61738 48685 61836 48706
rect 61738 48629 61759 48685
rect 61815 48629 61836 48685
rect 61738 48608 61836 48629
rect 63928 47944 64026 47961
rect 63928 47880 63945 47944
rect 64009 47880 64026 47944
rect 63928 47863 64026 47880
rect 1559 47336 1657 47353
rect 66163 47342 66261 47353
rect 1559 47272 1576 47336
rect 1640 47272 1657 47336
rect 1559 47255 1657 47272
rect 63939 47336 66261 47342
rect 63939 47272 63945 47336
rect 64009 47272 66180 47336
rect 66244 47272 66261 47336
rect 63939 47266 66261 47272
rect 66163 47255 66261 47266
rect 23962 46893 24060 46910
rect 23962 46829 23979 46893
rect 24043 46829 24060 46893
rect 23962 46812 24060 46829
rect 26458 46893 26556 46910
rect 26458 46829 26475 46893
rect 26539 46829 26556 46893
rect 26458 46812 26556 46829
rect 28954 46893 29052 46910
rect 28954 46829 28971 46893
rect 29035 46829 29052 46893
rect 28954 46812 29052 46829
rect 31450 46893 31548 46910
rect 31450 46829 31467 46893
rect 31531 46829 31548 46893
rect 31450 46812 31548 46829
rect 33946 46893 34044 46910
rect 33946 46829 33963 46893
rect 34027 46829 34044 46893
rect 33946 46812 34044 46829
rect 36442 46893 36540 46910
rect 36442 46829 36459 46893
rect 36523 46829 36540 46893
rect 36442 46812 36540 46829
rect 38938 46893 39036 46910
rect 38938 46829 38955 46893
rect 39019 46829 39036 46893
rect 38938 46812 39036 46829
rect 41434 46893 41532 46910
rect 41434 46829 41451 46893
rect 41515 46829 41532 46893
rect 41434 46812 41532 46829
rect 14130 46561 22074 46566
rect 14130 46560 41889 46561
rect 14130 46496 14136 46560
rect 14200 46496 22142 46560
rect 22206 46496 27297 46560
rect 27361 46496 40414 46560
rect 40478 46496 41889 46560
rect 14130 46495 41889 46496
rect 14130 46490 22074 46495
rect 21998 46238 41889 46239
rect 21998 46174 22004 46238
rect 22068 46174 41889 46238
rect 21998 46173 41889 46174
rect 1559 45656 1657 45673
rect 1559 45592 1576 45656
rect 1640 45592 1657 45656
rect 1559 45575 1657 45592
rect 66163 45656 66261 45673
rect 66163 45592 66180 45656
rect 66244 45592 66261 45656
rect 66163 45575 66261 45592
rect 21998 45400 41889 45401
rect 21998 45336 22004 45400
rect 22068 45336 41889 45400
rect 21998 45335 41889 45336
rect 21998 44626 41889 44627
rect 21998 44562 22142 44626
rect 22206 44562 41889 44626
rect 21998 44561 41889 44562
rect 46062 44391 46128 44394
rect 56951 44391 57017 44394
rect 46062 44389 57017 44391
rect 46062 44333 46067 44389
rect 46123 44333 56956 44389
rect 57012 44333 57017 44389
rect 46062 44331 57017 44333
rect 46062 44328 46128 44331
rect 56951 44328 57017 44331
rect 1559 43976 1657 43993
rect 66163 43982 66261 43993
rect 1559 43912 1576 43976
rect 1640 43912 1657 43976
rect 1559 43895 1657 43912
rect 64848 43976 66261 43982
rect 64848 43912 64854 43976
rect 64918 43912 66180 43976
rect 66244 43912 66261 43976
rect 64848 43906 66261 43912
rect 66163 43895 66261 43906
rect 46186 42993 46252 42996
rect 56951 42993 57017 42996
rect 46186 42991 57017 42993
rect 46186 42935 46191 42991
rect 46247 42935 56956 42991
rect 57012 42935 57017 42991
rect 46186 42933 57017 42935
rect 46186 42930 46252 42933
rect 56951 42930 57017 42933
rect 43199 42630 45324 42635
rect 21998 42629 45324 42630
rect 21998 42565 22142 42629
rect 22206 42565 22418 42629
rect 22482 42565 45254 42629
rect 45318 42565 45324 42629
rect 21998 42564 45324 42565
rect 43199 42559 45324 42564
rect 51639 42331 52296 42337
rect 1559 42302 1657 42313
rect 272 42296 1657 42302
rect 272 42232 278 42296
rect 342 42232 1576 42296
rect 1640 42232 1657 42296
rect 51639 42267 51645 42331
rect 51709 42267 52226 42331
rect 52290 42267 52296 42331
rect 66163 42302 66261 42313
rect 51639 42261 52296 42267
rect 64848 42296 67548 42302
rect 272 42226 1657 42232
rect 64848 42232 64854 42296
rect 64918 42292 67478 42296
rect 64918 42236 66184 42292
rect 66240 42236 67478 42292
rect 64918 42232 67478 42236
rect 67542 42232 67548 42296
rect 64848 42226 67548 42232
rect 1559 42215 1657 42226
rect 66163 42215 66261 42226
rect 65259 41846 65265 41848
rect 50344 41786 50404 41846
rect 56816 41786 65265 41846
rect 65259 41784 65265 41786
rect 65329 41784 65335 41848
rect 968 41619 10874 41625
rect 968 41555 974 41619
rect 1038 41555 10804 41619
rect 10868 41555 10874 41619
rect 968 41549 10874 41555
rect 49247 41579 49313 41582
rect 56951 41579 57017 41582
rect 49247 41577 57017 41579
rect 49247 41521 49252 41577
rect 49308 41521 56956 41577
rect 57012 41521 57017 41577
rect 49247 41519 57017 41521
rect 49247 41516 49313 41519
rect 56951 41516 57017 41519
rect 63744 41481 66852 41487
rect 63744 41417 63750 41481
rect 63814 41417 66782 41481
rect 66846 41417 66852 41481
rect 63744 41411 66852 41417
rect 44433 41097 45734 41102
rect 21998 41096 45734 41097
rect 21998 41032 22004 41096
rect 22068 41032 45664 41096
rect 45728 41032 45734 41096
rect 21998 41031 45734 41032
rect 44433 41026 45734 41031
rect 61830 41012 63820 41018
rect 61830 40948 61836 41012
rect 61900 40948 63750 41012
rect 63814 40948 63820 41012
rect 61830 40942 63820 40948
rect 1559 40616 1657 40633
rect 66163 40622 66261 40633
rect 1559 40552 1576 40616
rect 1640 40552 1657 40616
rect 1559 40535 1657 40552
rect 64848 40616 66261 40622
rect 64848 40552 64854 40616
rect 64918 40612 66261 40616
rect 64918 40556 66184 40612
rect 66240 40556 66261 40612
rect 64918 40552 66261 40556
rect 64848 40546 66261 40552
rect 66163 40535 66261 40546
rect 46748 40163 46846 40174
rect 45658 40157 46984 40163
rect 45658 40093 45664 40157
rect 45728 40093 46765 40157
rect 46829 40151 46984 40157
rect 48639 40151 48737 40162
rect 49471 40157 49569 40168
rect 48799 40151 50043 40157
rect 46829 40145 49973 40151
rect 46829 40093 48656 40145
rect 45658 40087 48656 40093
rect 46748 40076 46846 40087
rect 46908 40081 48656 40087
rect 48720 40087 49973 40145
rect 50037 40087 50043 40151
rect 48720 40081 50043 40087
rect 46908 40075 48875 40081
rect 48639 40064 48737 40075
rect 49471 40070 49569 40081
rect 1559 38936 1657 38953
rect 66163 38942 66261 38953
rect 1559 38872 1576 38936
rect 1640 38872 1657 38936
rect 1559 38855 1657 38872
rect 64848 38936 66261 38942
rect 64848 38872 64854 38936
rect 64918 38932 66261 38936
rect 64918 38876 66184 38932
rect 66240 38876 66261 38932
rect 64918 38872 66261 38876
rect 64848 38866 66261 38872
rect 66163 38855 66261 38866
rect 1559 37256 1657 37273
rect 66163 37262 66261 37273
rect 1559 37192 1576 37256
rect 1640 37192 1657 37256
rect 1559 37175 1657 37192
rect 66025 37252 66261 37262
rect 66025 37196 66184 37252
rect 66240 37196 66261 37252
rect 66025 37186 66261 37196
rect 66025 37169 66101 37186
rect 66163 37175 66261 37186
rect 64848 37163 66101 37169
rect 64848 37099 64854 37163
rect 64918 37099 66101 37163
rect 64848 37093 66101 37099
rect 1559 35576 1657 35593
rect 66163 35582 66261 35593
rect 1559 35512 1576 35576
rect 1640 35512 1657 35576
rect 1559 35495 1657 35512
rect 64848 35576 66261 35582
rect 64848 35512 64854 35576
rect 64918 35572 66261 35576
rect 64918 35516 66184 35572
rect 66240 35516 66261 35572
rect 64918 35512 66261 35516
rect 64848 35506 66261 35512
rect 66163 35495 66261 35506
rect 1559 33896 1657 33913
rect 66163 33902 66261 33913
rect 1559 33832 1576 33896
rect 1640 33832 1657 33896
rect 1559 33815 1657 33832
rect 64848 33896 66261 33902
rect 64848 33832 64854 33896
rect 64918 33892 66261 33896
rect 64918 33836 66184 33892
rect 66240 33836 66261 33892
rect 64918 33832 66261 33836
rect 64848 33826 66261 33832
rect 66163 33815 66261 33826
rect 1559 32222 1657 32233
rect 66163 32222 66261 32233
rect 272 32216 1657 32222
rect 272 32152 278 32216
rect 342 32152 1576 32216
rect 1640 32152 1657 32216
rect 272 32146 1657 32152
rect 64848 32216 67548 32222
rect 64848 32152 64854 32216
rect 64918 32212 67478 32216
rect 64918 32156 66184 32212
rect 66240 32156 67478 32212
rect 64918 32152 67478 32156
rect 67542 32152 67548 32216
rect 64848 32146 67548 32152
rect 1559 32135 1657 32146
rect 66163 32135 66261 32146
rect 65264 31645 65330 31646
rect 65222 31581 65265 31645
rect 65329 31581 65372 31645
rect 65264 31580 65330 31581
rect 968 31474 4076 31480
rect 968 31410 974 31474
rect 1038 31410 4006 31474
rect 4070 31410 4076 31474
rect 968 31404 4076 31410
rect 63744 31474 66852 31480
rect 63744 31410 63750 31474
rect 63814 31410 66782 31474
rect 66846 31410 66852 31474
rect 63744 31404 66852 31410
rect 1559 30542 1657 30553
rect 66163 30542 66261 30553
rect 272 30536 1657 30542
rect 272 30472 278 30536
rect 342 30472 1576 30536
rect 1640 30472 1657 30536
rect 272 30466 1657 30472
rect 64848 30536 66261 30542
rect 64848 30472 64854 30536
rect 64918 30472 66180 30536
rect 66244 30472 66261 30536
rect 64848 30466 66261 30472
rect 1559 30455 1657 30466
rect 66163 30455 66261 30466
rect 9789 30286 9887 30297
rect 0 30276 9887 30286
rect 0 30220 9810 30276
rect 9866 30220 9887 30276
rect 0 30210 9887 30220
rect 9789 30199 9887 30210
rect 10750 30207 10816 30210
rect 11404 30207 11470 30210
rect 10750 30205 11470 30207
rect 10750 30149 10755 30205
rect 10811 30149 11409 30205
rect 11465 30149 11470 30205
rect 10750 30147 11470 30149
rect 10750 30144 10816 30147
rect 11404 30144 11470 30147
rect 1559 28856 1657 28873
rect 1559 28792 1576 28856
rect 1640 28792 1657 28856
rect 1559 28775 1657 28792
rect 66163 28856 66261 28873
rect 66163 28792 66180 28856
rect 66244 28792 66261 28856
rect 66163 28775 66261 28792
rect 10750 28649 10816 28652
rect 11324 28649 11390 28652
rect 10750 28647 11390 28649
rect 9789 28586 9887 28597
rect 10750 28591 10755 28647
rect 10811 28591 11329 28647
rect 11385 28591 11390 28647
rect 10750 28589 11390 28591
rect 10750 28586 10816 28589
rect 11324 28586 11390 28589
rect 0 28576 9887 28586
rect 0 28520 9810 28576
rect 9866 28520 9887 28576
rect 0 28510 9887 28520
rect 9789 28499 9887 28510
rect 9789 27458 9887 27469
rect 0 27448 9887 27458
rect 0 27392 9810 27448
rect 9866 27392 9887 27448
rect 0 27382 9887 27392
rect 9789 27371 9887 27382
rect 10750 27379 10816 27382
rect 11244 27379 11310 27382
rect 10750 27377 11310 27379
rect 10750 27321 10755 27377
rect 10811 27321 11249 27377
rect 11305 27321 11310 27377
rect 10750 27319 11310 27321
rect 10750 27316 10816 27319
rect 11244 27316 11310 27319
rect 1559 27176 1657 27193
rect 1559 27112 1576 27176
rect 1640 27112 1657 27176
rect 1559 27095 1657 27112
rect 66163 27176 66261 27193
rect 66163 27112 66180 27176
rect 66244 27112 66261 27176
rect 66163 27095 66261 27112
rect 10750 25821 10816 25824
rect 11164 25821 11230 25824
rect 10750 25819 11230 25821
rect 9789 25758 9887 25769
rect 10750 25763 10755 25819
rect 10811 25763 11169 25819
rect 11225 25763 11230 25819
rect 10750 25761 11230 25763
rect 10750 25758 10816 25761
rect 11164 25758 11230 25761
rect 0 25748 9887 25758
rect 0 25692 9810 25748
rect 9866 25692 9887 25748
rect 0 25682 9887 25692
rect 9789 25671 9887 25682
rect 1559 25496 1657 25513
rect 1559 25432 1576 25496
rect 1640 25432 1657 25496
rect 1559 25415 1657 25432
rect 66163 25496 66261 25513
rect 66163 25432 66180 25496
rect 66244 25432 66261 25496
rect 66163 25415 66261 25432
rect 9789 24630 9887 24641
rect 0 24620 9887 24630
rect 0 24564 9810 24620
rect 9866 24564 9887 24620
rect 0 24554 9887 24564
rect 9789 24543 9887 24554
rect 10750 24551 10816 24554
rect 11084 24551 11150 24554
rect 10750 24549 11150 24551
rect 10750 24493 10755 24549
rect 10811 24493 11089 24549
rect 11145 24493 11150 24549
rect 10750 24491 11150 24493
rect 10750 24488 10816 24491
rect 11084 24488 11150 24491
rect 1559 23816 1657 23833
rect 1559 23752 1576 23816
rect 1640 23752 1657 23816
rect 1559 23735 1657 23752
rect 66163 23816 66261 23833
rect 66163 23752 66180 23816
rect 66244 23752 66261 23816
rect 66163 23735 66261 23752
rect 10750 22993 10816 22996
rect 11004 22993 11070 22996
rect 10750 22991 11070 22993
rect 9789 22930 9887 22941
rect 10750 22935 10755 22991
rect 10811 22935 11009 22991
rect 11065 22935 11070 22991
rect 10750 22933 11070 22935
rect 10750 22930 10816 22933
rect 11004 22930 11070 22933
rect 0 22920 9887 22930
rect 0 22864 9810 22920
rect 9866 22864 9887 22920
rect 0 22854 9887 22864
rect 9789 22843 9887 22854
rect 10836 22669 10920 22673
rect 10836 22664 10953 22669
rect 10836 22608 10892 22664
rect 10948 22608 10953 22664
rect 10836 22603 10953 22608
rect 10836 22599 10920 22603
rect 1719 22195 2972 22201
rect 1559 22142 1657 22153
rect 1719 22142 2902 22195
rect 1559 22136 2902 22142
rect 1559 22072 1576 22136
rect 1640 22131 2902 22136
rect 2966 22131 2972 22195
rect 1640 22125 2972 22131
rect 66163 22142 66261 22153
rect 66163 22136 67548 22142
rect 1640 22072 1795 22125
rect 1559 22066 1795 22072
rect 66163 22072 66180 22136
rect 66244 22072 67478 22136
rect 67542 22072 67548 22136
rect 66163 22066 67548 22072
rect 1559 22055 1657 22066
rect 66163 22055 66261 22066
rect 2490 21531 2556 21532
rect 2448 21467 2491 21531
rect 2555 21467 2598 21531
rect 2490 21466 2556 21467
rect 968 21328 4076 21334
rect 968 21264 974 21328
rect 1038 21264 4006 21328
rect 4070 21264 4076 21328
rect 968 21258 4076 21264
rect 63744 21328 66852 21334
rect 63744 21264 63750 21328
rect 63814 21264 66782 21328
rect 66846 21264 66852 21328
rect 63744 21258 66852 21264
rect 13960 20684 14581 20760
rect 13294 20612 13392 20629
rect 13294 20548 13311 20612
rect 13375 20548 13392 20612
rect 13294 20531 13392 20548
rect 13719 20618 13817 20629
rect 13960 20618 14036 20684
rect 14505 20622 14581 20684
rect 53402 20684 53857 20760
rect 13719 20612 14036 20618
rect 13719 20548 13736 20612
rect 13800 20548 14036 20612
rect 13719 20542 14036 20548
rect 14098 20611 14196 20622
rect 14098 20605 14432 20611
rect 13719 20531 13817 20542
rect 14098 20541 14115 20605
rect 14179 20541 14432 20605
rect 14098 20535 14432 20541
rect 14098 20524 14196 20535
rect 1559 20462 1657 20473
rect 272 20456 2972 20462
rect 272 20392 278 20456
rect 342 20452 2902 20456
rect 342 20396 1580 20452
rect 1636 20396 2902 20452
rect 342 20392 2902 20396
rect 2966 20392 2972 20456
rect 272 20386 2972 20392
rect 14356 20425 14432 20535
rect 14494 20524 14592 20622
rect 53144 20611 53242 20622
rect 53402 20611 53478 20684
rect 53144 20605 53478 20611
rect 53144 20541 53161 20605
rect 53225 20541 53478 20605
rect 53144 20535 53478 20541
rect 53540 20605 53638 20622
rect 53540 20541 53557 20605
rect 53621 20541 53638 20605
rect 53781 20618 53857 20684
rect 53919 20618 54017 20629
rect 53781 20542 54017 20618
rect 53144 20524 53242 20535
rect 53540 20524 53638 20541
rect 53919 20531 54017 20542
rect 54344 20612 54442 20629
rect 54344 20548 54361 20612
rect 54425 20548 54442 20612
rect 54344 20531 54442 20548
rect 66163 20462 66261 20473
rect 66163 20456 67548 20462
rect 14356 20419 16097 20425
rect 1559 20375 1657 20386
rect 14356 20355 16027 20419
rect 16091 20355 16097 20419
rect 66163 20392 66180 20456
rect 66244 20392 67478 20456
rect 67542 20392 67548 20456
rect 66163 20386 67548 20392
rect 66163 20375 66261 20386
rect 14356 20349 16097 20355
rect 9630 19964 12236 19970
rect 9630 19900 9636 19964
rect 9700 19900 12236 19964
rect 9630 19894 12236 19900
rect 12000 19821 12098 19832
rect 10798 19815 12098 19821
rect 10798 19751 10804 19815
rect 10868 19751 12017 19815
rect 12081 19751 12098 19815
rect 10798 19745 12098 19751
rect 12160 19821 12236 19894
rect 13960 19894 14581 19970
rect 12396 19821 12494 19832
rect 13294 19828 13392 19839
rect 13719 19828 13817 19839
rect 13960 19828 14036 19894
rect 14505 19832 14581 19894
rect 53155 19894 53776 19970
rect 53155 19832 53231 19894
rect 12694 19822 13392 19828
rect 12160 19745 12632 19821
rect 12694 19758 12700 19822
rect 12764 19758 13311 19822
rect 13375 19758 13392 19822
rect 12694 19752 13392 19758
rect 12000 19734 12098 19745
rect 12396 19734 12494 19745
rect 12556 19679 12632 19745
rect 13294 19741 13392 19752
rect 13454 19822 14036 19828
rect 13454 19758 13736 19822
rect 13800 19758 14036 19822
rect 13454 19752 14036 19758
rect 14098 19815 14196 19832
rect 13454 19679 13530 19752
rect 13719 19741 13817 19752
rect 14098 19751 14115 19815
rect 14179 19751 14196 19815
rect 14098 19734 14196 19751
rect 14494 19734 14592 19832
rect 53144 19815 53242 19832
rect 53144 19751 53161 19815
rect 53225 19751 53242 19815
rect 53144 19734 53242 19751
rect 53540 19815 53638 19832
rect 53540 19751 53557 19815
rect 53621 19751 53638 19815
rect 53700 19828 53776 19894
rect 54966 19894 55725 19970
rect 53919 19828 54017 19839
rect 54344 19828 54442 19839
rect 54966 19828 55042 19894
rect 55649 19832 55725 19894
rect 53700 19822 54282 19828
rect 53700 19758 53936 19822
rect 54000 19758 54282 19822
rect 53700 19752 54282 19758
rect 53540 19734 53638 19751
rect 53919 19741 54017 19752
rect 12556 19603 13530 19679
rect 54206 19679 54282 19752
rect 54344 19822 55042 19828
rect 54344 19758 54361 19822
rect 54425 19758 55042 19822
rect 55242 19821 55340 19832
rect 54344 19752 55042 19758
rect 54344 19741 54442 19752
rect 55104 19745 55340 19821
rect 55104 19679 55180 19745
rect 55242 19734 55340 19745
rect 55638 19734 55736 19832
rect 54206 19603 55180 19679
rect 12011 19535 12770 19541
rect 12011 19471 12017 19535
rect 12081 19471 12700 19535
rect 12764 19471 12770 19535
rect 12011 19465 12770 19471
rect 13305 19535 14185 19541
rect 13305 19471 13311 19535
rect 13375 19471 14115 19535
rect 14179 19471 14185 19535
rect 13305 19465 14185 19471
rect 53551 19535 54431 19541
rect 53551 19471 53557 19535
rect 53621 19471 54361 19535
rect 54425 19471 54431 19535
rect 53551 19465 54431 19471
rect 1719 18841 2972 18847
rect 1559 18782 1657 18793
rect 1719 18782 2902 18841
rect 1559 18777 2902 18782
rect 2966 18777 2972 18841
rect 1559 18772 2972 18777
rect 1559 18716 1580 18772
rect 1636 18771 2972 18772
rect 66163 18776 66261 18793
rect 1636 18716 1795 18771
rect 1559 18706 1795 18716
rect 66163 18712 66180 18776
rect 66244 18712 66261 18776
rect 1559 18695 1657 18706
rect 66163 18695 66261 18712
rect 13879 18314 14334 18390
rect 13294 18248 13392 18259
rect 13719 18248 13817 18259
rect 13879 18248 13955 18314
rect 13294 18242 13657 18248
rect 13294 18178 13311 18242
rect 13375 18178 13657 18242
rect 13294 18172 13657 18178
rect 13294 18161 13392 18172
rect 13581 18092 13657 18172
rect 13719 18242 13955 18248
rect 13719 18178 13736 18242
rect 13800 18178 13955 18242
rect 13719 18172 13955 18178
rect 14098 18235 14196 18252
rect 13719 18161 13817 18172
rect 14098 18171 14115 18235
rect 14179 18171 14196 18235
rect 14098 18154 14196 18171
rect 14258 18241 14334 18314
rect 53155 18314 53776 18390
rect 53155 18252 53231 18314
rect 14494 18241 14592 18252
rect 53144 18241 53242 18252
rect 14258 18235 14592 18241
rect 14258 18171 14511 18235
rect 14575 18171 14592 18235
rect 14258 18165 14592 18171
rect 51167 18235 53242 18241
rect 51167 18171 51173 18235
rect 51237 18171 53242 18235
rect 51167 18165 53242 18171
rect 14494 18154 14592 18165
rect 53144 18154 53242 18165
rect 53540 18235 53638 18252
rect 53540 18171 53557 18235
rect 53621 18171 53638 18235
rect 53700 18248 53776 18314
rect 53919 18248 54017 18259
rect 53700 18242 54017 18248
rect 53700 18178 53936 18242
rect 54000 18178 54017 18242
rect 53700 18172 54017 18178
rect 53540 18154 53638 18171
rect 53919 18161 54017 18172
rect 54344 18242 54442 18259
rect 54344 18178 54361 18242
rect 54425 18178 54442 18242
rect 54344 18161 54442 18178
rect 14109 18092 14185 18154
rect 13581 18016 14185 18092
rect 53551 17732 54431 17738
rect 53551 17668 53557 17732
rect 53621 17668 54361 17732
rect 54425 17668 54431 17732
rect 53551 17662 54431 17668
rect 12011 17524 12770 17600
rect 12011 17462 12087 17524
rect 12000 17364 12098 17462
rect 12396 17451 12494 17462
rect 12694 17458 12770 17524
rect 13879 17524 14334 17600
rect 13294 17458 13392 17469
rect 13719 17458 13817 17469
rect 13879 17458 13955 17524
rect 12694 17452 13392 17458
rect 12396 17375 12632 17451
rect 12694 17388 13311 17452
rect 13375 17388 13392 17452
rect 12694 17382 13392 17388
rect 12396 17364 12494 17375
rect 12556 17309 12632 17375
rect 13294 17371 13392 17382
rect 13454 17452 13955 17458
rect 13454 17388 13736 17452
rect 13800 17388 13955 17452
rect 13454 17382 13955 17388
rect 14098 17445 14196 17462
rect 13454 17309 13530 17382
rect 13719 17371 13817 17382
rect 14098 17381 14115 17445
rect 14179 17381 14196 17445
rect 14098 17364 14196 17381
rect 14258 17451 14334 17524
rect 53155 17524 53776 17600
rect 53155 17462 53231 17524
rect 14494 17451 14592 17462
rect 14258 17445 16569 17451
rect 14258 17381 14511 17445
rect 14575 17381 16499 17445
rect 16563 17381 16569 17445
rect 14258 17375 16569 17381
rect 14494 17364 14592 17375
rect 53144 17364 53242 17462
rect 53540 17445 53638 17462
rect 53540 17381 53557 17445
rect 53621 17381 53638 17445
rect 53700 17458 53776 17524
rect 54966 17524 55725 17600
rect 53919 17458 54017 17469
rect 54344 17458 54442 17469
rect 54966 17458 55042 17524
rect 55649 17462 55725 17524
rect 53700 17452 54282 17458
rect 53700 17388 53936 17452
rect 54000 17388 54282 17452
rect 53700 17382 54282 17388
rect 53540 17364 53638 17381
rect 53919 17371 54017 17382
rect 12556 17233 13530 17309
rect 53551 17265 53627 17364
rect 51639 17259 53627 17265
rect 51639 17195 51645 17259
rect 51709 17195 53627 17259
rect 54206 17309 54282 17382
rect 54344 17452 55042 17458
rect 54344 17388 54361 17452
rect 54425 17388 55042 17452
rect 55242 17451 55340 17462
rect 54344 17382 55042 17388
rect 54344 17371 54442 17382
rect 55104 17375 55340 17451
rect 55104 17309 55180 17375
rect 55242 17364 55340 17375
rect 55638 17364 55736 17462
rect 54206 17233 55180 17309
rect 51639 17189 53627 17195
rect 1559 17102 1657 17113
rect 1559 17092 1795 17102
rect 1559 17036 1580 17092
rect 1636 17081 1795 17092
rect 66163 17096 66261 17113
rect 1636 17075 2972 17081
rect 1636 17036 2902 17075
rect 1559 17026 2902 17036
rect 1559 17015 1657 17026
rect 1719 17011 2902 17026
rect 2966 17011 2972 17075
rect 66163 17032 66180 17096
rect 66244 17032 66261 17096
rect 66163 17015 66261 17032
rect 1719 17005 2972 17011
rect 13960 15944 14581 16020
rect 13294 15878 13392 15889
rect 13719 15878 13817 15889
rect 13960 15878 14036 15944
rect 14505 15882 14581 15944
rect 53402 15944 53857 16020
rect 13294 15872 13657 15878
rect 13294 15808 13311 15872
rect 13375 15808 13657 15872
rect 13294 15802 13657 15808
rect 13294 15791 13392 15802
rect 13581 15722 13657 15802
rect 13719 15872 14036 15878
rect 13719 15808 13736 15872
rect 13800 15808 14036 15872
rect 13719 15802 14036 15808
rect 14098 15865 14196 15882
rect 13719 15791 13817 15802
rect 14098 15801 14115 15865
rect 14179 15801 14196 15865
rect 14098 15784 14196 15801
rect 14494 15865 14592 15882
rect 14494 15801 14511 15865
rect 14575 15801 14592 15865
rect 14494 15784 14592 15801
rect 53144 15871 53242 15882
rect 53402 15871 53478 15944
rect 53144 15865 53478 15871
rect 53144 15801 53161 15865
rect 53225 15801 53478 15865
rect 53144 15795 53478 15801
rect 53540 15865 53638 15882
rect 53540 15801 53557 15865
rect 53621 15801 53638 15865
rect 53781 15878 53857 15944
rect 53919 15878 54017 15889
rect 54344 15878 54442 15889
rect 53781 15872 54017 15878
rect 53781 15808 53936 15872
rect 54000 15808 54017 15872
rect 53781 15802 54017 15808
rect 53144 15784 53242 15795
rect 53540 15784 53638 15801
rect 53919 15791 54017 15802
rect 54079 15872 54442 15878
rect 54079 15808 54361 15872
rect 54425 15808 54442 15872
rect 54079 15802 54442 15808
rect 14109 15722 14185 15784
rect 13581 15646 14185 15722
rect 53551 15722 53627 15784
rect 54079 15722 54155 15802
rect 54344 15791 54442 15802
rect 53551 15646 54155 15722
rect 19653 15470 22488 15476
rect 1559 15422 1657 15433
rect 1559 15416 2972 15422
rect 1559 15412 2902 15416
rect 1559 15356 1580 15412
rect 1636 15356 2902 15412
rect 1559 15352 2902 15356
rect 2966 15352 2972 15416
rect 19653 15406 19659 15470
rect 19723 15406 22418 15470
rect 22482 15406 22488 15470
rect 19653 15400 22488 15406
rect 66163 15416 66261 15433
rect 1559 15346 2972 15352
rect 66163 15352 66180 15416
rect 66244 15352 66261 15416
rect 1559 15335 1657 15346
rect 66163 15335 66261 15352
rect 12011 15154 12770 15230
rect 12011 15092 12087 15154
rect 12000 15081 12098 15092
rect 12396 15081 12494 15092
rect 12694 15088 12770 15154
rect 13879 15154 14334 15230
rect 13294 15088 13392 15099
rect 13719 15088 13817 15099
rect 13879 15088 13955 15154
rect 12694 15082 13392 15088
rect 5914 15075 12098 15081
rect 5914 15011 5920 15075
rect 5984 15011 12098 15075
rect 5914 15005 12098 15011
rect 12000 14994 12098 15005
rect 12160 15005 12632 15081
rect 12694 15018 13311 15082
rect 13375 15018 13392 15082
rect 12694 15012 13392 15018
rect 12160 14932 12236 15005
rect 12396 14994 12494 15005
rect 10714 14926 12236 14932
rect 10714 14862 10720 14926
rect 10784 14862 12236 14926
rect 12556 14939 12632 15005
rect 13294 15001 13392 15012
rect 13454 15012 13955 15088
rect 14098 15075 14196 15092
rect 13454 14939 13530 15012
rect 13719 15001 13817 15012
rect 14098 15011 14115 15075
rect 14179 15011 14196 15075
rect 14098 14994 14196 15011
rect 14258 15081 14334 15154
rect 53155 15154 53776 15230
rect 53155 15092 53231 15154
rect 14494 15081 14592 15092
rect 14258 15075 14592 15081
rect 14258 15011 14511 15075
rect 14575 15011 14592 15075
rect 53144 15075 53242 15092
rect 45248 15055 51715 15061
rect 14258 15005 14592 15011
rect 14494 14994 14592 15005
rect 16021 15027 19729 15033
rect 16021 14963 16027 15027
rect 16091 14963 17275 15027
rect 17339 14963 18591 15027
rect 18655 14963 19659 15027
rect 19723 14963 19729 15027
rect 45248 14991 45254 15055
rect 45318 14991 48013 15055
rect 48077 14991 49081 15055
rect 49145 14991 50397 15055
rect 50461 14991 51645 15055
rect 51709 14991 51715 15055
rect 53144 15011 53161 15075
rect 53225 15011 53242 15075
rect 53144 14994 53242 15011
rect 53540 15075 53638 15092
rect 53540 15011 53557 15075
rect 53621 15011 53638 15075
rect 53700 15088 53776 15154
rect 54355 15161 55725 15237
rect 54355 15099 54431 15161
rect 53919 15088 54017 15099
rect 53700 15012 54017 15088
rect 53540 14994 53638 15011
rect 53919 15001 54017 15012
rect 54344 15082 54442 15099
rect 55649 15092 55725 15161
rect 54344 15018 54361 15082
rect 54425 15018 54442 15082
rect 55242 15081 55340 15092
rect 54344 15001 54442 15018
rect 54504 15005 55340 15081
rect 45248 14985 51715 14991
rect 16021 14957 19729 14963
rect 12556 14863 13530 14939
rect 53930 14939 54006 15001
rect 54504 14939 54580 15005
rect 55242 14994 55340 15005
rect 55638 15081 55736 15092
rect 55638 15075 57022 15081
rect 55638 15011 56952 15075
rect 57016 15011 57022 15075
rect 55638 15005 57022 15011
rect 55638 14994 55736 15005
rect 53930 14863 54580 14939
rect 55253 14932 55329 14994
rect 55253 14926 58190 14932
rect 10714 14856 12236 14862
rect 55253 14862 58120 14926
rect 58184 14862 58190 14926
rect 55253 14856 58190 14862
rect 16493 14685 17769 14691
rect 16493 14621 16499 14685
rect 16563 14621 16931 14685
rect 16995 14621 17699 14685
rect 17763 14621 17769 14685
rect 16493 14615 17769 14621
rect 49967 14685 51243 14691
rect 49967 14621 49973 14685
rect 50037 14621 50741 14685
rect 50805 14621 51173 14685
rect 51237 14621 51243 14685
rect 49967 14615 51243 14621
rect 18167 14495 18265 14506
rect 18999 14501 19097 14512
rect 18327 14495 19235 14501
rect 17693 14489 19016 14495
rect 17693 14425 17699 14489
rect 17763 14431 19016 14489
rect 19080 14489 19235 14495
rect 20890 14489 20988 14500
rect 19080 14483 22078 14489
rect 19080 14431 20907 14483
rect 17763 14425 20907 14431
rect 17693 14419 18403 14425
rect 18167 14408 18265 14419
rect 18999 14414 19097 14425
rect 19159 14419 20907 14425
rect 20971 14419 22008 14483
rect 22072 14419 22078 14483
rect 19159 14413 22078 14419
rect 20890 14402 20988 14413
rect 56900 14373 56984 14377
rect 56867 14368 56984 14373
rect 56867 14312 56872 14368
rect 56928 14312 56984 14368
rect 56867 14307 56984 14312
rect 56900 14303 56984 14307
rect 57933 14122 58031 14133
rect 57933 14112 67820 14122
rect 57933 14056 57954 14112
rect 58010 14056 67820 14112
rect 57933 14046 67820 14056
rect 56666 14043 56732 14046
rect 57004 14043 57070 14046
rect 56666 14041 57070 14043
rect 56666 13985 56671 14041
rect 56727 13985 57009 14041
rect 57065 13985 57070 14041
rect 57933 14035 58031 14046
rect 56666 13983 57070 13985
rect 56666 13980 56732 13983
rect 57004 13980 57070 13983
rect 1559 13742 1657 13753
rect 1559 13736 2972 13742
rect 1559 13732 2902 13736
rect 1559 13676 1580 13732
rect 1636 13676 2902 13732
rect 1559 13672 2902 13676
rect 2966 13672 2972 13736
rect 1559 13666 2972 13672
rect 66163 13736 66261 13753
rect 66163 13672 66180 13736
rect 66244 13672 66261 13736
rect 1559 13655 1657 13666
rect 66163 13655 66261 13672
rect 21998 13494 43885 13495
rect 21998 13430 22004 13494
rect 22068 13430 23634 13494
rect 23698 13430 43885 13494
rect 21998 13429 43885 13430
rect 10803 13007 10869 13010
rect 18423 13007 18489 13010
rect 10803 13005 18489 13007
rect 10803 12949 10808 13005
rect 10864 12949 18428 13005
rect 18484 12949 18489 13005
rect 10803 12947 18489 12949
rect 10803 12944 10869 12947
rect 18423 12944 18489 12947
rect 2485 12678 2491 12742
rect 2555 12740 2561 12742
rect 2555 12680 23804 12740
rect 2555 12678 2561 12680
rect 56586 12485 56652 12488
rect 57004 12485 57070 12488
rect 56586 12483 57070 12485
rect 56586 12427 56591 12483
rect 56647 12427 57009 12483
rect 57065 12427 57070 12483
rect 56586 12425 57070 12427
rect 56586 12422 56652 12425
rect 57004 12422 57070 12425
rect 57933 12422 58031 12433
rect 57933 12412 67820 12422
rect 57933 12356 57954 12412
rect 58010 12356 67820 12412
rect 57933 12346 67820 12356
rect 57933 12335 58031 12346
rect 15440 12259 16097 12265
rect 15440 12195 15446 12259
rect 15510 12195 16027 12259
rect 16091 12195 16097 12259
rect 15440 12189 16097 12195
rect 1559 12062 1657 12073
rect 1559 12056 2972 12062
rect 1559 12052 2902 12056
rect 1559 11996 1580 12052
rect 1636 11996 2902 12052
rect 1559 11992 2902 11996
rect 2966 11992 2972 12056
rect 1559 11986 2972 11992
rect 66163 12056 66261 12073
rect 66163 11992 66180 12056
rect 66244 11992 66261 12056
rect 1559 11975 1657 11986
rect 66163 11975 66261 11992
rect 21998 11961 43275 11962
rect 21998 11897 22004 11961
rect 22068 11897 22418 11961
rect 22482 11897 43275 11961
rect 21998 11896 43275 11897
rect 57933 11294 58031 11305
rect 57933 11284 67820 11294
rect 57933 11228 57954 11284
rect 58010 11228 67820 11284
rect 57933 11218 67820 11228
rect 56506 11215 56572 11218
rect 57004 11215 57070 11218
rect 56506 11213 57070 11215
rect 968 11183 4076 11189
rect 968 11119 974 11183
rect 1038 11119 4006 11183
rect 4070 11119 4076 11183
rect 56506 11157 56511 11213
rect 56567 11157 57009 11213
rect 57065 11157 57070 11213
rect 57933 11207 58031 11218
rect 56506 11155 57070 11157
rect 56506 11152 56572 11155
rect 57004 11152 57070 11155
rect 968 11113 4076 11119
rect 56946 11079 66852 11085
rect 56946 11015 56952 11079
rect 57016 11015 66782 11079
rect 66846 11015 66852 11079
rect 56946 11009 66852 11015
rect 1559 10382 1657 10393
rect 66163 10382 66261 10393
rect 272 10376 2972 10382
rect 272 10312 278 10376
rect 342 10372 2902 10376
rect 342 10316 1580 10372
rect 1636 10316 2902 10372
rect 342 10312 2902 10316
rect 2966 10312 2972 10376
rect 272 10306 2972 10312
rect 66163 10376 67548 10382
rect 66163 10312 66180 10376
rect 66244 10312 67478 10376
rect 67542 10312 67548 10376
rect 66163 10306 67548 10312
rect 1559 10295 1657 10306
rect 66163 10295 66261 10306
rect 10803 10179 10869 10182
rect 21450 10179 21516 10182
rect 10803 10177 21516 10179
rect 10803 10121 10808 10177
rect 10864 10121 21455 10177
rect 21511 10121 21516 10177
rect 10803 10119 21516 10121
rect 10803 10116 10869 10119
rect 21450 10116 21516 10119
rect 21998 9745 41889 9746
rect 21998 9681 22004 9745
rect 22068 9681 23496 9745
rect 23560 9681 41889 9745
rect 21998 9680 41889 9681
rect 56426 9657 56492 9660
rect 57004 9657 57070 9660
rect 56426 9655 57070 9657
rect 4000 9612 5990 9618
rect 4000 9548 4006 9612
rect 4070 9548 5920 9612
rect 5984 9548 5990 9612
rect 56426 9599 56431 9655
rect 56487 9599 57009 9655
rect 57065 9599 57070 9655
rect 56426 9597 57070 9599
rect 56426 9594 56492 9597
rect 57004 9594 57070 9597
rect 57933 9594 58031 9605
rect 4000 9542 5990 9548
rect 57657 9588 58031 9594
rect 57657 9524 57663 9588
rect 57727 9584 58031 9588
rect 57727 9528 57954 9584
rect 58010 9528 58031 9584
rect 57727 9524 58031 9528
rect 57657 9518 58031 9524
rect 57933 9507 58031 9518
rect 21998 9308 41889 9309
rect 21998 9244 22004 9308
rect 22068 9244 23634 9308
rect 23698 9244 41889 9308
rect 21998 9243 41889 9244
rect 21998 8976 41889 8977
rect 21998 8912 23496 8976
rect 23560 8912 40414 8976
rect 40478 8912 41889 8976
rect 21998 8911 41889 8912
rect 10803 8765 10869 8768
rect 21574 8765 21640 8768
rect 10803 8763 21640 8765
rect 1559 8702 1657 8713
rect 10803 8707 10808 8763
rect 10864 8707 21579 8763
rect 21635 8707 21640 8763
rect 10803 8705 21640 8707
rect 10803 8702 10869 8705
rect 21574 8702 21640 8705
rect 1559 8696 2972 8702
rect 1559 8632 1576 8696
rect 1640 8632 2902 8696
rect 2966 8632 2972 8696
rect 1559 8626 2972 8632
rect 66163 8696 66261 8713
rect 66163 8632 66180 8696
rect 66244 8632 66261 8696
rect 1559 8615 1657 8626
rect 66163 8615 66261 8632
rect 21998 8484 41889 8485
rect 21998 8420 22004 8484
rect 22068 8420 41889 8484
rect 57933 8466 58031 8477
rect 21998 8419 41889 8420
rect 57795 8460 58031 8466
rect 57795 8396 57801 8460
rect 57865 8456 58031 8460
rect 57865 8400 57954 8456
rect 58010 8400 58031 8456
rect 57865 8396 58031 8400
rect 57795 8390 58031 8396
rect 56346 8387 56412 8390
rect 57004 8387 57070 8390
rect 56346 8385 57070 8387
rect 56346 8329 56351 8385
rect 56407 8329 57009 8385
rect 57065 8329 57070 8385
rect 57933 8379 58031 8390
rect 56346 8327 57070 8329
rect 56346 8324 56412 8327
rect 57004 8324 57070 8327
rect 1559 7016 1657 7033
rect 1559 6952 1576 7016
rect 1640 6952 1657 7016
rect 1559 6935 1657 6952
rect 66163 7016 66261 7033
rect 66163 6952 66180 7016
rect 66244 6952 66261 7016
rect 66163 6935 66261 6952
rect 56266 6829 56332 6832
rect 57004 6829 57070 6832
rect 56266 6827 57070 6829
rect 56266 6771 56271 6827
rect 56327 6771 57009 6827
rect 57065 6771 57070 6827
rect 56266 6769 57070 6771
rect 56266 6766 56332 6769
rect 57004 6766 57070 6769
rect 57933 6760 58031 6777
rect 57933 6696 57950 6760
rect 58014 6696 58031 6760
rect 57933 6679 58031 6696
rect 1559 5342 1657 5353
rect 1559 5336 3732 5342
rect 1559 5272 1576 5336
rect 1640 5272 3732 5336
rect 1559 5266 3732 5272
rect 1559 5255 1657 5266
rect 3656 5238 3732 5266
rect 66163 5336 66261 5353
rect 66163 5272 66180 5336
rect 66244 5272 66261 5336
rect 66163 5255 66261 5272
rect 3794 5238 3892 5249
rect 3656 5162 3892 5238
rect 3794 5151 3892 5162
rect 5984 4483 6082 4504
rect 5984 4427 6005 4483
rect 6061 4427 6082 4483
rect 5984 4406 6082 4427
rect 2687 4388 2785 4399
rect 0 4378 2785 4388
rect 0 4322 2708 4378
rect 2764 4322 2785 4378
rect 0 4312 2785 4322
rect 2687 4301 2785 4312
rect 5995 4344 6071 4406
rect 5995 4338 6128 4344
rect 5995 4274 6058 4338
rect 6122 4274 6128 4338
rect 5995 4268 6128 4274
rect 11955 3900 12053 3911
rect 10714 3894 12053 3900
rect 3794 3824 3892 3835
rect 10714 3830 10720 3894
rect 10784 3830 11972 3894
rect 12036 3830 12053 3894
rect 10714 3824 12053 3830
rect 3794 3818 5809 3824
rect 3794 3754 5739 3818
rect 5803 3754 5809 3818
rect 11955 3813 12053 3824
rect 14291 3894 14389 3911
rect 18963 3900 19061 3911
rect 14291 3830 14308 3894
rect 14372 3830 14389 3894
rect 14291 3813 14389 3830
rect 18706 3894 19061 3900
rect 18706 3830 18712 3894
rect 18776 3830 19061 3894
rect 18706 3824 19061 3830
rect 18963 3813 19061 3824
rect 3794 3748 5809 3754
rect 3794 3737 3892 3748
rect 1559 3656 1657 3673
rect 1559 3592 1576 3656
rect 1640 3592 1657 3656
rect 1559 3575 1657 3592
rect 66163 3656 66261 3673
rect 66163 3592 66180 3656
rect 66244 3592 66261 3656
rect 66163 3575 66261 3592
rect 12125 3044 12223 3061
rect 12125 2980 12142 3044
rect 12206 2980 12223 3044
rect 12125 2963 12223 2980
rect 13293 3044 13391 3061
rect 13293 2980 13310 3044
rect 13374 2980 13391 3044
rect 13293 2963 13391 2980
rect 14461 3044 14559 3061
rect 14461 2980 14478 3044
rect 14542 2980 14559 3044
rect 14461 2963 14559 2980
rect 15629 3044 15727 3061
rect 15629 2980 15646 3044
rect 15710 2980 15727 3044
rect 15629 2963 15727 2980
rect 16797 3044 16895 3061
rect 16797 2980 16814 3044
rect 16878 2980 16895 3044
rect 16797 2963 16895 2980
rect 17965 3044 18063 3061
rect 17965 2980 17982 3044
rect 18046 2980 18063 3044
rect 17965 2963 18063 2980
rect 19133 3044 19231 3061
rect 19133 2980 19150 3044
rect 19214 2980 19231 3044
rect 19133 2963 19231 2980
rect 20301 3044 20399 3061
rect 20301 2980 20318 3044
rect 20382 2980 20399 3044
rect 20301 2963 20399 2980
rect 21469 3044 21567 3061
rect 21469 2980 21486 3044
rect 21550 2980 21567 3044
rect 21469 2963 21567 2980
rect 22637 3044 22735 3061
rect 22637 2980 22654 3044
rect 22718 2980 22735 3044
rect 22637 2963 22735 2980
rect 10887 2786 10953 2789
rect 10887 2784 13172 2786
rect 10887 2728 10892 2784
rect 10948 2728 13172 2784
rect 10887 2726 13172 2728
rect 10887 2723 10953 2726
rect 13123 2480 13221 2497
rect 15459 2486 15557 2497
rect 20131 2486 20229 2497
rect 13123 2416 13140 2480
rect 13204 2416 13221 2480
rect 13123 2399 13221 2416
rect 14130 2480 27367 2486
rect 14130 2416 14136 2480
rect 14200 2416 15285 2480
rect 15349 2416 27297 2480
rect 27361 2416 27367 2480
rect 14130 2410 27367 2416
rect 15459 2399 15557 2410
rect 20131 2399 20229 2410
rect 1559 1976 1657 1993
rect 66163 1982 66261 1993
rect 1559 1912 1576 1976
rect 1640 1912 1657 1976
rect 1559 1895 1657 1912
rect 65746 1976 66261 1982
rect 65746 1912 65752 1976
rect 65816 1912 66180 1976
rect 66244 1912 66261 1976
rect 65746 1906 66261 1912
rect 66163 1895 66261 1906
rect 1895 1646 1993 1657
rect 3575 1646 3673 1657
rect 5255 1646 5353 1657
rect 6935 1646 7033 1657
rect 8615 1646 8713 1657
rect 10295 1646 10393 1657
rect 11975 1646 12073 1657
rect 13655 1646 13753 1657
rect 15335 1646 15433 1657
rect 17015 1646 17113 1657
rect 18695 1646 18793 1657
rect 20375 1646 20473 1657
rect 22055 1646 22153 1657
rect 23735 1646 23833 1657
rect 25415 1646 25513 1657
rect 27095 1646 27193 1657
rect 28775 1646 28873 1657
rect 30455 1646 30553 1657
rect 32135 1646 32233 1657
rect 33815 1646 33913 1657
rect 35495 1646 35593 1657
rect 37175 1646 37273 1657
rect 38855 1646 38953 1657
rect 40535 1646 40633 1657
rect 42215 1646 42313 1657
rect 43895 1646 43993 1657
rect 45575 1646 45673 1657
rect 47255 1646 47353 1657
rect 48935 1646 49033 1657
rect 50615 1646 50713 1657
rect 52295 1646 52393 1657
rect 53975 1646 54073 1657
rect 55655 1646 55753 1657
rect 57335 1646 57433 1657
rect 59015 1646 59113 1657
rect 60695 1646 60793 1657
rect 1570 1640 60793 1646
rect 1570 1576 1576 1640
rect 1640 1636 11992 1640
rect 1640 1580 1916 1636
rect 1972 1580 3596 1636
rect 3652 1580 5276 1636
rect 5332 1580 6956 1636
rect 7012 1580 8636 1636
rect 8692 1580 10316 1636
rect 10372 1580 11992 1636
rect 1640 1576 11992 1580
rect 12056 1576 13672 1640
rect 13736 1576 14308 1640
rect 14372 1636 18712 1640
rect 18776 1636 27112 1640
rect 27176 1636 40552 1640
rect 40616 1636 53992 1640
rect 54056 1636 60793 1640
rect 14372 1580 15356 1636
rect 15412 1580 17036 1636
rect 17092 1580 18712 1636
rect 18776 1580 20396 1636
rect 20452 1580 22076 1636
rect 22132 1580 23756 1636
rect 23812 1580 25436 1636
rect 25492 1580 27112 1636
rect 27176 1580 28796 1636
rect 28852 1580 30476 1636
rect 30532 1580 32156 1636
rect 32212 1580 33836 1636
rect 33892 1580 35516 1636
rect 35572 1580 37196 1636
rect 37252 1580 38876 1636
rect 38932 1580 40552 1636
rect 40616 1580 42236 1636
rect 42292 1580 43916 1636
rect 43972 1580 45596 1636
rect 45652 1580 47276 1636
rect 47332 1580 48956 1636
rect 49012 1580 50636 1636
rect 50692 1580 52316 1636
rect 52372 1580 53992 1636
rect 54056 1580 55676 1636
rect 55732 1580 57356 1636
rect 57412 1580 59036 1636
rect 59092 1580 60716 1636
rect 60772 1580 60793 1636
rect 14372 1576 18712 1580
rect 18776 1576 27112 1580
rect 27176 1576 40552 1580
rect 40616 1576 53992 1580
rect 54056 1576 60793 1580
rect 1570 1570 60793 1576
rect 1895 1559 1993 1570
rect 3575 1559 3673 1570
rect 5255 1559 5353 1570
rect 6935 1559 7033 1570
rect 8615 1559 8713 1570
rect 10295 1559 10393 1570
rect 11975 1559 12073 1570
rect 13655 1559 13753 1570
rect 15335 1559 15433 1570
rect 17015 1559 17113 1570
rect 18695 1559 18793 1570
rect 20375 1559 20473 1570
rect 22055 1559 22153 1570
rect 23735 1559 23833 1570
rect 25415 1559 25513 1570
rect 27095 1559 27193 1570
rect 28775 1559 28873 1570
rect 30455 1559 30553 1570
rect 32135 1559 32233 1570
rect 33815 1559 33913 1570
rect 35495 1559 35593 1570
rect 37175 1559 37273 1570
rect 38855 1559 38953 1570
rect 40535 1559 40633 1570
rect 42215 1559 42313 1570
rect 43895 1559 43993 1570
rect 45575 1559 45673 1570
rect 47255 1559 47353 1570
rect 48935 1559 49033 1570
rect 50615 1559 50713 1570
rect 52295 1559 52393 1570
rect 53975 1559 54073 1570
rect 55655 1559 55753 1570
rect 57335 1559 57433 1570
rect 59015 1559 59113 1570
rect 60695 1559 60793 1570
rect 62375 1646 62473 1657
rect 64055 1646 64153 1657
rect 65735 1646 65833 1657
rect 62375 1640 65833 1646
rect 62375 1636 65752 1640
rect 62375 1580 62396 1636
rect 62452 1580 64076 1636
rect 64132 1580 65752 1636
rect 62375 1576 65752 1580
rect 65816 1576 65833 1640
rect 62375 1570 65833 1576
rect 62375 1559 62473 1570
rect 64055 1559 64153 1570
rect 65735 1559 65833 1570
rect 696 1038 67124 1044
rect 696 974 702 1038
rect 766 974 838 1038
rect 902 974 974 1038
rect 1038 974 13140 1038
rect 13204 974 14136 1038
rect 14200 974 27297 1038
rect 27361 974 40414 1038
rect 40478 974 56952 1038
rect 57016 974 66782 1038
rect 66846 974 66918 1038
rect 66982 974 67054 1038
rect 67118 974 67124 1038
rect 696 902 67124 974
rect 696 838 702 902
rect 766 838 838 902
rect 902 838 974 902
rect 1038 838 66782 902
rect 66846 838 66918 902
rect 66982 838 67054 902
rect 67118 838 67124 902
rect 696 766 67124 838
rect 696 702 702 766
rect 766 702 838 766
rect 902 702 974 766
rect 1038 702 66782 766
rect 66846 702 66918 766
rect 66982 702 67054 766
rect 67118 702 67124 766
rect 696 696 67124 702
rect 0 342 67820 348
rect 0 278 6 342
rect 70 278 142 342
rect 206 278 278 342
rect 342 278 13672 342
rect 13736 278 27112 342
rect 27176 278 40552 342
rect 40616 278 53992 342
rect 54056 278 67478 342
rect 67542 278 67614 342
rect 67678 278 67750 342
rect 67814 278 67820 342
rect 0 206 67820 278
rect 0 142 6 206
rect 70 142 142 206
rect 206 142 278 206
rect 342 142 67478 206
rect 67542 142 67614 206
rect 67678 142 67750 206
rect 67814 142 67820 206
rect 0 70 67820 142
rect 0 6 6 70
rect 70 6 142 70
rect 206 6 278 70
rect 342 6 67478 70
rect 67542 6 67614 70
rect 67678 6 67750 70
rect 67814 6 67820 70
rect 0 0 67820 6
<< via3 >>
rect 6 52668 70 52732
rect 142 52668 206 52732
rect 278 52668 342 52732
rect 67478 52668 67542 52732
rect 67614 52668 67678 52732
rect 67750 52668 67814 52732
rect 6 52532 70 52596
rect 142 52532 206 52596
rect 278 52532 342 52596
rect 67478 52532 67542 52596
rect 67614 52532 67678 52596
rect 67750 52532 67814 52596
rect 6 52396 70 52460
rect 142 52396 206 52460
rect 278 52396 342 52460
rect 13672 52396 13736 52460
rect 27112 52396 27176 52460
rect 40552 52396 40616 52460
rect 53992 52396 54056 52460
rect 67478 52396 67542 52460
rect 67614 52396 67678 52460
rect 67750 52396 67814 52460
rect 702 51972 766 52036
rect 838 51972 902 52036
rect 974 51972 1038 52036
rect 66782 51972 66846 52036
rect 66918 51972 66982 52036
rect 67054 51972 67118 52036
rect 702 51836 766 51900
rect 838 51836 902 51900
rect 974 51836 1038 51900
rect 66782 51836 66846 51900
rect 66918 51836 66982 51900
rect 67054 51836 67118 51900
rect 702 51700 766 51764
rect 838 51700 902 51764
rect 974 51700 1038 51764
rect 14136 51700 14200 51764
rect 27297 51700 27361 51764
rect 40414 51700 40478 51764
rect 53448 51700 53512 51764
rect 66782 51700 66846 51764
rect 66918 51700 66982 51764
rect 67054 51700 67118 51764
rect 1912 51158 1976 51162
rect 13672 51158 13736 51162
rect 27112 51158 27176 51162
rect 40552 51158 40616 51162
rect 53992 51158 54056 51162
rect 1912 51102 1916 51158
rect 1916 51102 1972 51158
rect 1972 51102 1976 51158
rect 13672 51102 13676 51158
rect 13676 51102 13732 51158
rect 13732 51102 13736 51158
rect 27112 51102 27116 51158
rect 27116 51102 27172 51158
rect 27172 51102 27176 51158
rect 40552 51102 40556 51158
rect 40556 51102 40612 51158
rect 40612 51102 40616 51158
rect 53992 51102 53996 51158
rect 53996 51102 54052 51158
rect 54052 51102 54056 51158
rect 1912 51098 1976 51102
rect 13672 51098 13736 51102
rect 27112 51098 27176 51102
rect 40552 51098 40616 51102
rect 53992 51098 54056 51102
rect 54616 51098 54680 51162
rect 66180 51098 66244 51162
rect 1576 50692 1640 50696
rect 1576 50636 1580 50692
rect 1580 50636 1636 50692
rect 1636 50636 1640 50692
rect 1576 50632 1640 50636
rect 1912 50632 1976 50696
rect 66180 50692 66244 50696
rect 66180 50636 66184 50692
rect 66184 50636 66240 50692
rect 66240 50636 66244 50692
rect 66180 50632 66244 50636
rect 52226 50258 52290 50322
rect 53448 50258 53512 50322
rect 61836 50258 61900 50322
rect 53278 49754 53342 49758
rect 53278 49698 53282 49754
rect 53282 49698 53338 49754
rect 53338 49698 53342 49754
rect 53278 49694 53342 49698
rect 54446 49754 54510 49758
rect 54446 49698 54450 49754
rect 54450 49698 54506 49754
rect 54506 49698 54510 49754
rect 54446 49694 54510 49698
rect 62017 49294 62081 49358
rect 1576 49012 1640 49016
rect 1576 48956 1580 49012
rect 1580 48956 1636 49012
rect 1636 48956 1640 49012
rect 1576 48952 1640 48956
rect 66180 49012 66244 49016
rect 66180 48956 66184 49012
rect 66184 48956 66240 49012
rect 66240 48956 66244 49012
rect 66180 48952 66244 48956
rect 54616 48844 54680 48908
rect 57036 48844 57100 48908
rect 61698 48774 61762 48838
rect 63945 47880 64009 47944
rect 1576 47332 1640 47336
rect 1576 47276 1580 47332
rect 1580 47276 1636 47332
rect 1636 47276 1640 47332
rect 1576 47272 1640 47276
rect 63945 47272 64009 47336
rect 66180 47332 66244 47336
rect 66180 47276 66184 47332
rect 66184 47276 66240 47332
rect 66240 47276 66244 47332
rect 66180 47272 66244 47276
rect 23979 46889 24043 46893
rect 23979 46833 23983 46889
rect 23983 46833 24039 46889
rect 24039 46833 24043 46889
rect 23979 46829 24043 46833
rect 26475 46889 26539 46893
rect 26475 46833 26479 46889
rect 26479 46833 26535 46889
rect 26535 46833 26539 46889
rect 26475 46829 26539 46833
rect 28971 46889 29035 46893
rect 28971 46833 28975 46889
rect 28975 46833 29031 46889
rect 29031 46833 29035 46889
rect 28971 46829 29035 46833
rect 31467 46889 31531 46893
rect 31467 46833 31471 46889
rect 31471 46833 31527 46889
rect 31527 46833 31531 46889
rect 31467 46829 31531 46833
rect 33963 46889 34027 46893
rect 33963 46833 33967 46889
rect 33967 46833 34023 46889
rect 34023 46833 34027 46889
rect 33963 46829 34027 46833
rect 36459 46889 36523 46893
rect 36459 46833 36463 46889
rect 36463 46833 36519 46889
rect 36519 46833 36523 46889
rect 36459 46829 36523 46833
rect 38955 46889 39019 46893
rect 38955 46833 38959 46889
rect 38959 46833 39015 46889
rect 39015 46833 39019 46889
rect 38955 46829 39019 46833
rect 41451 46889 41515 46893
rect 41451 46833 41455 46889
rect 41455 46833 41511 46889
rect 41511 46833 41515 46889
rect 41451 46829 41515 46833
rect 14136 46496 14200 46560
rect 22142 46496 22206 46560
rect 27297 46496 27361 46560
rect 40414 46496 40478 46560
rect 22004 46174 22068 46238
rect 1576 45652 1640 45656
rect 1576 45596 1580 45652
rect 1580 45596 1636 45652
rect 1636 45596 1640 45652
rect 1576 45592 1640 45596
rect 66180 45652 66244 45656
rect 66180 45596 66184 45652
rect 66184 45596 66240 45652
rect 66240 45596 66244 45652
rect 66180 45592 66244 45596
rect 22004 45336 22068 45400
rect 22142 44562 22206 44626
rect 1576 43972 1640 43976
rect 1576 43916 1580 43972
rect 1580 43916 1636 43972
rect 1636 43916 1640 43972
rect 1576 43912 1640 43916
rect 64854 43912 64918 43976
rect 66180 43972 66244 43976
rect 66180 43916 66184 43972
rect 66184 43916 66240 43972
rect 66240 43916 66244 43972
rect 66180 43912 66244 43916
rect 22142 42565 22206 42629
rect 22418 42565 22482 42629
rect 45254 42565 45318 42629
rect 278 42232 342 42296
rect 1576 42292 1640 42296
rect 1576 42236 1580 42292
rect 1580 42236 1636 42292
rect 1636 42236 1640 42292
rect 1576 42232 1640 42236
rect 51645 42267 51709 42331
rect 52226 42267 52290 42331
rect 64854 42232 64918 42296
rect 67478 42232 67542 42296
rect 65265 41784 65329 41848
rect 974 41555 1038 41619
rect 10804 41555 10868 41619
rect 63750 41417 63814 41481
rect 66782 41417 66846 41481
rect 22004 41032 22068 41096
rect 45664 41032 45728 41096
rect 61836 40948 61900 41012
rect 63750 40948 63814 41012
rect 1576 40612 1640 40616
rect 1576 40556 1580 40612
rect 1580 40556 1636 40612
rect 1636 40556 1640 40612
rect 1576 40552 1640 40556
rect 64854 40552 64918 40616
rect 45664 40093 45728 40157
rect 46765 40153 46829 40157
rect 46765 40097 46769 40153
rect 46769 40097 46825 40153
rect 46825 40097 46829 40153
rect 46765 40093 46829 40097
rect 48656 40141 48720 40145
rect 48656 40085 48660 40141
rect 48660 40085 48716 40141
rect 48716 40085 48720 40141
rect 49973 40087 50037 40151
rect 48656 40081 48720 40085
rect 1576 38932 1640 38936
rect 1576 38876 1580 38932
rect 1580 38876 1636 38932
rect 1636 38876 1640 38932
rect 1576 38872 1640 38876
rect 64854 38872 64918 38936
rect 1576 37252 1640 37256
rect 1576 37196 1580 37252
rect 1580 37196 1636 37252
rect 1636 37196 1640 37252
rect 1576 37192 1640 37196
rect 64854 37099 64918 37163
rect 1576 35572 1640 35576
rect 1576 35516 1580 35572
rect 1580 35516 1636 35572
rect 1636 35516 1640 35572
rect 1576 35512 1640 35516
rect 64854 35512 64918 35576
rect 1576 33892 1640 33896
rect 1576 33836 1580 33892
rect 1580 33836 1636 33892
rect 1636 33836 1640 33892
rect 1576 33832 1640 33836
rect 64854 33832 64918 33896
rect 278 32152 342 32216
rect 1576 32212 1640 32216
rect 1576 32156 1580 32212
rect 1580 32156 1636 32212
rect 1636 32156 1640 32212
rect 1576 32152 1640 32156
rect 64854 32152 64918 32216
rect 67478 32152 67542 32216
rect 65265 31641 65329 31645
rect 65265 31585 65269 31641
rect 65269 31585 65325 31641
rect 65325 31585 65329 31641
rect 65265 31581 65329 31585
rect 974 31410 1038 31474
rect 4006 31410 4070 31474
rect 63750 31410 63814 31474
rect 66782 31410 66846 31474
rect 278 30472 342 30536
rect 1576 30532 1640 30536
rect 1576 30476 1580 30532
rect 1580 30476 1636 30532
rect 1636 30476 1640 30532
rect 1576 30472 1640 30476
rect 64854 30472 64918 30536
rect 66180 30532 66244 30536
rect 66180 30476 66184 30532
rect 66184 30476 66240 30532
rect 66240 30476 66244 30532
rect 66180 30472 66244 30476
rect 1576 28852 1640 28856
rect 1576 28796 1580 28852
rect 1580 28796 1636 28852
rect 1636 28796 1640 28852
rect 1576 28792 1640 28796
rect 66180 28852 66244 28856
rect 66180 28796 66184 28852
rect 66184 28796 66240 28852
rect 66240 28796 66244 28852
rect 66180 28792 66244 28796
rect 1576 27172 1640 27176
rect 1576 27116 1580 27172
rect 1580 27116 1636 27172
rect 1636 27116 1640 27172
rect 1576 27112 1640 27116
rect 66180 27172 66244 27176
rect 66180 27116 66184 27172
rect 66184 27116 66240 27172
rect 66240 27116 66244 27172
rect 66180 27112 66244 27116
rect 1576 25492 1640 25496
rect 1576 25436 1580 25492
rect 1580 25436 1636 25492
rect 1636 25436 1640 25492
rect 1576 25432 1640 25436
rect 66180 25492 66244 25496
rect 66180 25436 66184 25492
rect 66184 25436 66240 25492
rect 66240 25436 66244 25492
rect 66180 25432 66244 25436
rect 1576 23812 1640 23816
rect 1576 23756 1580 23812
rect 1580 23756 1636 23812
rect 1636 23756 1640 23812
rect 1576 23752 1640 23756
rect 66180 23812 66244 23816
rect 66180 23756 66184 23812
rect 66184 23756 66240 23812
rect 66240 23756 66244 23812
rect 66180 23752 66244 23756
rect 1576 22132 1640 22136
rect 1576 22076 1580 22132
rect 1580 22076 1636 22132
rect 1636 22076 1640 22132
rect 2902 22131 2966 22195
rect 1576 22072 1640 22076
rect 66180 22132 66244 22136
rect 66180 22076 66184 22132
rect 66184 22076 66240 22132
rect 66240 22076 66244 22132
rect 66180 22072 66244 22076
rect 67478 22072 67542 22136
rect 2491 21527 2555 21531
rect 2491 21471 2495 21527
rect 2495 21471 2551 21527
rect 2551 21471 2555 21527
rect 2491 21467 2555 21471
rect 974 21264 1038 21328
rect 4006 21264 4070 21328
rect 63750 21264 63814 21328
rect 66782 21264 66846 21328
rect 13311 20548 13375 20612
rect 13736 20548 13800 20612
rect 14115 20541 14179 20605
rect 278 20392 342 20456
rect 2902 20392 2966 20456
rect 53161 20541 53225 20605
rect 53557 20541 53621 20605
rect 54361 20548 54425 20612
rect 16027 20355 16091 20419
rect 66180 20452 66244 20456
rect 66180 20396 66184 20452
rect 66184 20396 66240 20452
rect 66240 20396 66244 20452
rect 66180 20392 66244 20396
rect 67478 20392 67542 20456
rect 9636 19900 9700 19964
rect 10804 19751 10868 19815
rect 12017 19751 12081 19815
rect 12700 19758 12764 19822
rect 13311 19758 13375 19822
rect 13736 19758 13800 19822
rect 14115 19751 14179 19815
rect 53161 19751 53225 19815
rect 53557 19751 53621 19815
rect 53936 19758 54000 19822
rect 54361 19758 54425 19822
rect 12017 19471 12081 19535
rect 12700 19471 12764 19535
rect 13311 19471 13375 19535
rect 14115 19471 14179 19535
rect 53557 19471 53621 19535
rect 54361 19471 54425 19535
rect 2902 18777 2966 18841
rect 66180 18772 66244 18776
rect 66180 18716 66184 18772
rect 66184 18716 66240 18772
rect 66240 18716 66244 18772
rect 66180 18712 66244 18716
rect 13311 18178 13375 18242
rect 13736 18178 13800 18242
rect 14115 18171 14179 18235
rect 14511 18171 14575 18235
rect 51173 18171 51237 18235
rect 53557 18171 53621 18235
rect 53936 18178 54000 18242
rect 54361 18178 54425 18242
rect 53557 17668 53621 17732
rect 54361 17668 54425 17732
rect 13311 17388 13375 17452
rect 13736 17388 13800 17452
rect 14115 17381 14179 17445
rect 14511 17381 14575 17445
rect 16499 17381 16563 17445
rect 53557 17381 53621 17445
rect 53936 17388 54000 17452
rect 51645 17195 51709 17259
rect 54361 17388 54425 17452
rect 2902 17011 2966 17075
rect 66180 17092 66244 17096
rect 66180 17036 66184 17092
rect 66184 17036 66240 17092
rect 66240 17036 66244 17092
rect 66180 17032 66244 17036
rect 13311 15808 13375 15872
rect 13736 15808 13800 15872
rect 14115 15801 14179 15865
rect 14511 15801 14575 15865
rect 53161 15801 53225 15865
rect 53557 15801 53621 15865
rect 53936 15808 54000 15872
rect 54361 15808 54425 15872
rect 2902 15352 2966 15416
rect 19659 15406 19723 15470
rect 22418 15406 22482 15470
rect 66180 15412 66244 15416
rect 66180 15356 66184 15412
rect 66184 15356 66240 15412
rect 66240 15356 66244 15412
rect 66180 15352 66244 15356
rect 5920 15011 5984 15075
rect 13311 15018 13375 15082
rect 10720 14862 10784 14926
rect 14115 15011 14179 15075
rect 14511 15011 14575 15075
rect 16027 14963 16091 15027
rect 17275 14963 17339 15027
rect 18591 14963 18655 15027
rect 19659 14963 19723 15027
rect 45254 14991 45318 15055
rect 48013 14991 48077 15055
rect 49081 14991 49145 15055
rect 50397 14991 50461 15055
rect 51645 14991 51709 15055
rect 53161 15011 53225 15075
rect 53557 15011 53621 15075
rect 54361 15018 54425 15082
rect 56952 15011 57016 15075
rect 58120 14862 58184 14926
rect 16499 14621 16563 14685
rect 16931 14621 16995 14685
rect 17699 14621 17763 14685
rect 49973 14621 50037 14685
rect 50741 14621 50805 14685
rect 51173 14621 51237 14685
rect 19016 14491 19080 14495
rect 17699 14425 17763 14489
rect 19016 14435 19020 14491
rect 19020 14435 19076 14491
rect 19076 14435 19080 14491
rect 19016 14431 19080 14435
rect 20907 14479 20971 14483
rect 20907 14423 20911 14479
rect 20911 14423 20967 14479
rect 20967 14423 20971 14479
rect 20907 14419 20971 14423
rect 22008 14419 22072 14483
rect 2902 13672 2966 13736
rect 66180 13732 66244 13736
rect 66180 13676 66184 13732
rect 66184 13676 66240 13732
rect 66240 13676 66244 13732
rect 66180 13672 66244 13676
rect 22004 13430 22068 13494
rect 23634 13430 23698 13494
rect 2491 12678 2555 12742
rect 15446 12195 15510 12259
rect 16027 12195 16091 12259
rect 2902 11992 2966 12056
rect 66180 12052 66244 12056
rect 66180 11996 66184 12052
rect 66184 11996 66240 12052
rect 66240 11996 66244 12052
rect 66180 11992 66244 11996
rect 22004 11897 22068 11961
rect 22418 11897 22482 11961
rect 974 11119 1038 11183
rect 4006 11119 4070 11183
rect 56952 11015 57016 11079
rect 66782 11015 66846 11079
rect 278 10312 342 10376
rect 2902 10312 2966 10376
rect 66180 10372 66244 10376
rect 66180 10316 66184 10372
rect 66184 10316 66240 10372
rect 66240 10316 66244 10372
rect 66180 10312 66244 10316
rect 67478 10312 67542 10376
rect 22004 9681 22068 9745
rect 23496 9681 23560 9745
rect 4006 9548 4070 9612
rect 5920 9548 5984 9612
rect 57663 9524 57727 9588
rect 22004 9244 22068 9308
rect 23634 9244 23698 9308
rect 23496 8912 23560 8976
rect 40414 8912 40478 8976
rect 1576 8692 1640 8696
rect 1576 8636 1580 8692
rect 1580 8636 1636 8692
rect 1636 8636 1640 8692
rect 1576 8632 1640 8636
rect 2902 8632 2966 8696
rect 66180 8692 66244 8696
rect 66180 8636 66184 8692
rect 66184 8636 66240 8692
rect 66240 8636 66244 8692
rect 66180 8632 66244 8636
rect 22004 8420 22068 8484
rect 57801 8396 57865 8460
rect 1576 7012 1640 7016
rect 1576 6956 1580 7012
rect 1580 6956 1636 7012
rect 1636 6956 1640 7012
rect 1576 6952 1640 6956
rect 66180 7012 66244 7016
rect 66180 6956 66184 7012
rect 66184 6956 66240 7012
rect 66240 6956 66244 7012
rect 66180 6952 66244 6956
rect 57950 6756 58014 6760
rect 57950 6700 57954 6756
rect 57954 6700 58010 6756
rect 58010 6700 58014 6756
rect 57950 6696 58014 6700
rect 1576 5332 1640 5336
rect 1576 5276 1580 5332
rect 1580 5276 1636 5332
rect 1636 5276 1640 5332
rect 1576 5272 1640 5276
rect 66180 5332 66244 5336
rect 66180 5276 66184 5332
rect 66184 5276 66240 5332
rect 66240 5276 66244 5332
rect 66180 5272 66244 5276
rect 6058 4274 6122 4338
rect 10720 3830 10784 3894
rect 11972 3830 12036 3894
rect 5739 3754 5803 3818
rect 14308 3830 14372 3894
rect 18712 3830 18776 3894
rect 1576 3652 1640 3656
rect 1576 3596 1580 3652
rect 1580 3596 1636 3652
rect 1636 3596 1640 3652
rect 1576 3592 1640 3596
rect 66180 3652 66244 3656
rect 66180 3596 66184 3652
rect 66184 3596 66240 3652
rect 66240 3596 66244 3652
rect 66180 3592 66244 3596
rect 12142 3040 12206 3044
rect 12142 2984 12146 3040
rect 12146 2984 12202 3040
rect 12202 2984 12206 3040
rect 12142 2980 12206 2984
rect 13310 3040 13374 3044
rect 13310 2984 13314 3040
rect 13314 2984 13370 3040
rect 13370 2984 13374 3040
rect 13310 2980 13374 2984
rect 14478 3040 14542 3044
rect 14478 2984 14482 3040
rect 14482 2984 14538 3040
rect 14538 2984 14542 3040
rect 14478 2980 14542 2984
rect 15646 3040 15710 3044
rect 15646 2984 15650 3040
rect 15650 2984 15706 3040
rect 15706 2984 15710 3040
rect 15646 2980 15710 2984
rect 16814 3040 16878 3044
rect 16814 2984 16818 3040
rect 16818 2984 16874 3040
rect 16874 2984 16878 3040
rect 16814 2980 16878 2984
rect 17982 3040 18046 3044
rect 17982 2984 17986 3040
rect 17986 2984 18042 3040
rect 18042 2984 18046 3040
rect 17982 2980 18046 2984
rect 19150 3040 19214 3044
rect 19150 2984 19154 3040
rect 19154 2984 19210 3040
rect 19210 2984 19214 3040
rect 19150 2980 19214 2984
rect 20318 3040 20382 3044
rect 20318 2984 20322 3040
rect 20322 2984 20378 3040
rect 20378 2984 20382 3040
rect 20318 2980 20382 2984
rect 21486 3040 21550 3044
rect 21486 2984 21490 3040
rect 21490 2984 21546 3040
rect 21546 2984 21550 3040
rect 21486 2980 21550 2984
rect 22654 3040 22718 3044
rect 22654 2984 22658 3040
rect 22658 2984 22714 3040
rect 22714 2984 22718 3040
rect 22654 2980 22718 2984
rect 13140 2416 13204 2480
rect 14136 2416 14200 2480
rect 15285 2416 15349 2480
rect 27297 2416 27361 2480
rect 1576 1972 1640 1976
rect 1576 1916 1580 1972
rect 1580 1916 1636 1972
rect 1636 1916 1640 1972
rect 1576 1912 1640 1916
rect 65752 1912 65816 1976
rect 66180 1972 66244 1976
rect 66180 1916 66184 1972
rect 66184 1916 66240 1972
rect 66240 1916 66244 1972
rect 66180 1912 66244 1916
rect 1576 1576 1640 1640
rect 11992 1636 12056 1640
rect 11992 1580 11996 1636
rect 11996 1580 12052 1636
rect 12052 1580 12056 1636
rect 11992 1576 12056 1580
rect 13672 1636 13736 1640
rect 13672 1580 13676 1636
rect 13676 1580 13732 1636
rect 13732 1580 13736 1636
rect 13672 1576 13736 1580
rect 14308 1576 14372 1640
rect 18712 1636 18776 1640
rect 27112 1636 27176 1640
rect 40552 1636 40616 1640
rect 53992 1636 54056 1640
rect 18712 1580 18716 1636
rect 18716 1580 18772 1636
rect 18772 1580 18776 1636
rect 27112 1580 27116 1636
rect 27116 1580 27172 1636
rect 27172 1580 27176 1636
rect 40552 1580 40556 1636
rect 40556 1580 40612 1636
rect 40612 1580 40616 1636
rect 53992 1580 53996 1636
rect 53996 1580 54052 1636
rect 54052 1580 54056 1636
rect 18712 1576 18776 1580
rect 27112 1576 27176 1580
rect 40552 1576 40616 1580
rect 53992 1576 54056 1580
rect 65752 1636 65816 1640
rect 65752 1580 65756 1636
rect 65756 1580 65812 1636
rect 65812 1580 65816 1636
rect 65752 1576 65816 1580
rect 702 974 766 1038
rect 838 974 902 1038
rect 974 974 1038 1038
rect 13140 974 13204 1038
rect 14136 974 14200 1038
rect 27297 974 27361 1038
rect 40414 974 40478 1038
rect 56952 974 57016 1038
rect 66782 974 66846 1038
rect 66918 974 66982 1038
rect 67054 974 67118 1038
rect 702 838 766 902
rect 838 838 902 902
rect 974 838 1038 902
rect 66782 838 66846 902
rect 66918 838 66982 902
rect 67054 838 67118 902
rect 702 702 766 766
rect 838 702 902 766
rect 974 702 1038 766
rect 66782 702 66846 766
rect 66918 702 66982 766
rect 67054 702 67118 766
rect 6 278 70 342
rect 142 278 206 342
rect 278 278 342 342
rect 13672 278 13736 342
rect 27112 278 27176 342
rect 40552 278 40616 342
rect 53992 278 54056 342
rect 67478 278 67542 342
rect 67614 278 67678 342
rect 67750 278 67814 342
rect 6 142 70 206
rect 142 142 206 206
rect 278 142 342 206
rect 67478 142 67542 206
rect 67614 142 67678 206
rect 67750 142 67814 206
rect 6 6 70 70
rect 142 6 206 70
rect 278 6 342 70
rect 67478 6 67542 70
rect 67614 6 67678 70
rect 67750 6 67814 70
<< metal4 >>
rect 0 52732 348 52738
rect 0 52668 6 52732
rect 70 52668 142 52732
rect 206 52668 278 52732
rect 342 52668 348 52732
rect 0 52596 348 52668
rect 0 52532 6 52596
rect 70 52532 142 52596
rect 206 52532 278 52596
rect 342 52532 348 52596
rect 0 52460 348 52532
rect 0 52396 6 52460
rect 70 52396 142 52460
rect 206 52396 278 52460
rect 342 52396 348 52460
rect 0 42296 348 52396
rect 13666 52460 13742 52466
rect 13666 52396 13672 52460
rect 13736 52396 13742 52460
rect 0 42232 278 42296
rect 342 42232 348 42296
rect 0 32216 348 42232
rect 0 32152 278 32216
rect 342 32152 348 32216
rect 0 30536 348 32152
rect 0 30472 278 30536
rect 342 30472 348 30536
rect 0 20456 348 30472
rect 0 20392 278 20456
rect 342 20392 348 20456
rect 0 10376 348 20392
rect 0 10312 278 10376
rect 342 10312 348 10376
rect 0 342 348 10312
rect 696 52036 1044 52042
rect 696 51972 702 52036
rect 766 51972 838 52036
rect 902 51972 974 52036
rect 1038 51972 1044 52036
rect 696 51900 1044 51972
rect 696 51836 702 51900
rect 766 51836 838 51900
rect 902 51836 974 51900
rect 1038 51836 1044 51900
rect 696 51764 1044 51836
rect 696 51700 702 51764
rect 766 51700 838 51764
rect 902 51700 974 51764
rect 1038 51700 1044 51764
rect 696 41619 1044 51700
rect 1906 51162 1982 51168
rect 1906 51098 1912 51162
rect 1976 51098 1982 51162
rect 696 41555 974 41619
rect 1038 41555 1044 41619
rect 696 31474 1044 41555
rect 1570 50696 1646 50702
rect 1570 50632 1576 50696
rect 1640 50632 1646 50696
rect 1570 49016 1646 50632
rect 1906 50696 1982 51098
rect 13666 51162 13742 52396
rect 13666 51098 13672 51162
rect 13736 51098 13742 51162
rect 13666 51092 13742 51098
rect 14130 51764 14206 51770
rect 14130 51700 14136 51764
rect 14200 51700 14206 51764
rect 1906 50632 1912 50696
rect 1976 50632 1982 50696
rect 1906 50626 1982 50632
rect 1570 48952 1576 49016
rect 1640 48952 1646 49016
rect 1570 47336 1646 48952
rect 1570 47272 1576 47336
rect 1640 47272 1646 47336
rect 1570 45656 1646 47272
rect 14130 46560 14206 51700
rect 23973 46893 24049 52738
rect 23973 46829 23979 46893
rect 24043 46829 24049 46893
rect 23973 46823 24049 46829
rect 26469 46893 26545 52738
rect 27106 52460 27182 52466
rect 27106 52396 27112 52460
rect 27176 52396 27182 52460
rect 27106 51162 27182 52396
rect 27106 51098 27112 51162
rect 27176 51098 27182 51162
rect 27106 51092 27182 51098
rect 27291 51764 27367 51770
rect 27291 51700 27297 51764
rect 27361 51700 27367 51764
rect 26469 46829 26475 46893
rect 26539 46829 26545 46893
rect 26469 46823 26545 46829
rect 14130 46496 14136 46560
rect 14200 46496 14206 46560
rect 14130 46490 14206 46496
rect 22136 46560 22212 46566
rect 22136 46496 22142 46560
rect 22206 46496 22212 46560
rect 1570 45592 1576 45656
rect 1640 45592 1646 45656
rect 1570 43976 1646 45592
rect 1570 43912 1576 43976
rect 1640 43912 1646 43976
rect 1570 42296 1646 43912
rect 1570 42232 1576 42296
rect 1640 42232 1646 42296
rect 1570 40616 1646 42232
rect 21998 46238 22074 46244
rect 21998 46174 22004 46238
rect 22068 46174 22074 46238
rect 21998 45400 22074 46174
rect 21998 45336 22004 45400
rect 22068 45336 22074 45400
rect 1570 40552 1576 40616
rect 1640 40552 1646 40616
rect 1570 38936 1646 40552
rect 1570 38872 1576 38936
rect 1640 38872 1646 38936
rect 1570 37256 1646 38872
rect 1570 37192 1576 37256
rect 1640 37192 1646 37256
rect 1570 35576 1646 37192
rect 1570 35512 1576 35576
rect 1640 35512 1646 35576
rect 1570 33896 1646 35512
rect 1570 33832 1576 33896
rect 1640 33832 1646 33896
rect 1570 32216 1646 33832
rect 1570 32152 1576 32216
rect 1640 32152 1646 32216
rect 1570 32146 1646 32152
rect 10798 41619 10874 41625
rect 10798 41555 10804 41619
rect 10868 41555 10874 41619
rect 696 31410 974 31474
rect 1038 31410 1044 31474
rect 696 21328 1044 31410
rect 4000 31474 4076 31480
rect 4000 31410 4006 31474
rect 4070 31410 4076 31474
rect 1570 30536 1646 30542
rect 1570 30472 1576 30536
rect 1640 30472 1646 30536
rect 1570 28856 1646 30472
rect 1570 28792 1576 28856
rect 1640 28792 1646 28856
rect 1570 27176 1646 28792
rect 1570 27112 1576 27176
rect 1640 27112 1646 27176
rect 1570 25496 1646 27112
rect 1570 25432 1576 25496
rect 1640 25432 1646 25496
rect 1570 23816 1646 25432
rect 1570 23752 1576 23816
rect 1640 23752 1646 23816
rect 1570 22136 1646 23752
rect 1570 22072 1576 22136
rect 1640 22072 1646 22136
rect 1570 22066 1646 22072
rect 2901 22195 2967 22201
rect 2901 22131 2902 22195
rect 2966 22131 2967 22195
rect 4000 22142 4076 31410
rect 9635 22371 9701 30845
rect 10798 30787 10874 41555
rect 21998 41096 22074 45336
rect 22136 44626 22212 46496
rect 27291 46560 27367 51700
rect 28965 46893 29041 52738
rect 28965 46829 28971 46893
rect 29035 46829 29041 46893
rect 28965 46823 29041 46829
rect 31461 46893 31537 52738
rect 31461 46829 31467 46893
rect 31531 46829 31537 46893
rect 31461 46823 31537 46829
rect 33957 46893 34033 52738
rect 33957 46829 33963 46893
rect 34027 46829 34033 46893
rect 33957 46823 34033 46829
rect 36453 46893 36529 52738
rect 36453 46829 36459 46893
rect 36523 46829 36529 46893
rect 36453 46823 36529 46829
rect 38949 46893 39025 52738
rect 40546 52460 40622 52466
rect 40546 52396 40552 52460
rect 40616 52396 40622 52460
rect 38949 46829 38955 46893
rect 39019 46829 39025 46893
rect 38949 46823 39025 46829
rect 40408 51764 40484 51770
rect 40408 51700 40414 51764
rect 40478 51700 40484 51764
rect 27291 46496 27297 46560
rect 27361 46496 27367 46560
rect 27291 46490 27367 46496
rect 40408 46560 40484 51700
rect 40546 51162 40622 52396
rect 40546 51098 40552 51162
rect 40616 51098 40622 51162
rect 40546 51092 40622 51098
rect 41445 46893 41521 52738
rect 52220 50322 52296 50328
rect 52220 50258 52226 50322
rect 52290 50258 52296 50322
rect 41445 46829 41451 46893
rect 41515 46829 41521 46893
rect 41445 46823 41521 46829
rect 40408 46496 40414 46560
rect 40478 46496 40484 46560
rect 40408 46490 40484 46496
rect 22136 44562 22142 44626
rect 22206 44562 22212 44626
rect 22136 42629 22212 44562
rect 22136 42565 22142 42629
rect 22206 42565 22212 42629
rect 22136 42559 22212 42565
rect 22412 42629 22488 42635
rect 22412 42565 22418 42629
rect 22482 42565 22488 42629
rect 21998 41032 22004 41096
rect 22068 41032 22074 41096
rect 21998 40861 22074 41032
rect 21998 40785 22078 40861
rect 22002 40642 22078 40785
rect 22412 40642 22488 42565
rect 45248 42629 45324 42635
rect 45248 42565 45254 42629
rect 45318 42565 45324 42629
rect 45248 40642 45324 42565
rect 51015 42529 51081 48175
rect 52220 48148 52296 50258
rect 53272 49758 53348 52738
rect 53986 52460 54062 52466
rect 53986 52396 53992 52460
rect 54056 52396 54062 52460
rect 53442 51764 53518 51770
rect 53442 51700 53448 51764
rect 53512 51700 53518 51764
rect 53442 50322 53518 51700
rect 53986 51162 54062 52396
rect 53986 51098 53992 51162
rect 54056 51098 54062 51162
rect 53986 51092 54062 51098
rect 53442 50258 53448 50322
rect 53512 50258 53518 50322
rect 53442 50252 53518 50258
rect 53272 49694 53278 49758
rect 53342 49694 53348 49758
rect 53272 49688 53348 49694
rect 54440 49758 54516 52738
rect 54440 49694 54446 49758
rect 54510 49694 54516 49758
rect 54440 49688 54516 49694
rect 54610 51162 54686 51168
rect 54610 51098 54616 51162
rect 54680 51098 54686 51162
rect 54610 48908 54686 51098
rect 54610 48844 54616 48908
rect 54680 48844 54686 48908
rect 54610 48838 54686 48844
rect 57030 48908 57106 48914
rect 57030 48844 57036 48908
rect 57100 48844 57106 48908
rect 51010 42453 51243 42529
rect 52225 42480 52291 48148
rect 57030 47869 57106 48844
rect 61692 48838 61768 52738
rect 67472 52732 67820 52738
rect 67472 52668 67478 52732
rect 67542 52668 67614 52732
rect 67678 52668 67750 52732
rect 67814 52668 67820 52732
rect 67472 52596 67820 52668
rect 67472 52532 67478 52596
rect 67542 52532 67614 52596
rect 67678 52532 67750 52596
rect 67814 52532 67820 52596
rect 67472 52460 67820 52532
rect 67472 52396 67478 52460
rect 67542 52396 67614 52460
rect 67678 52396 67750 52460
rect 67814 52396 67820 52460
rect 66776 52036 67124 52042
rect 66776 51972 66782 52036
rect 66846 51972 66918 52036
rect 66982 51972 67054 52036
rect 67118 51972 67124 52036
rect 66776 51900 67124 51972
rect 66776 51836 66782 51900
rect 66846 51836 66918 51900
rect 66982 51836 67054 51900
rect 67118 51836 67124 51900
rect 66776 51764 67124 51836
rect 66776 51700 66782 51764
rect 66846 51700 66918 51764
rect 66982 51700 67054 51764
rect 67118 51700 67124 51764
rect 66174 51162 66250 51168
rect 66174 51098 66180 51162
rect 66244 51098 66250 51162
rect 66174 50696 66250 51098
rect 66174 50632 66180 50696
rect 66244 50632 66250 50696
rect 61830 50322 61906 50328
rect 61830 50258 61836 50322
rect 61900 50258 61906 50322
rect 61830 49359 61906 50258
rect 62011 49359 62087 49364
rect 61830 49358 62087 49359
rect 61830 49294 62017 49358
rect 62081 49294 62087 49358
rect 61830 49283 62087 49294
rect 61692 48774 61698 48838
rect 61762 48774 61768 48838
rect 61692 48768 61768 48774
rect 45658 41096 45734 41102
rect 45658 41032 45664 41096
rect 45728 41032 45734 41096
rect 45658 40642 45734 41032
rect 2490 21531 2556 21532
rect 2490 21467 2491 21531
rect 2555 21467 2556 21531
rect 2490 21466 2556 21467
rect 696 21264 974 21328
rect 1038 21264 1044 21328
rect 696 11183 1044 21264
rect 2493 12743 2553 21466
rect 2901 20456 2967 22131
rect 2901 20392 2902 20456
rect 2966 20392 2967 20456
rect 2901 18841 2967 20392
rect 2901 18777 2902 18841
rect 2966 18777 2967 18841
rect 2901 17075 2967 18777
rect 2901 17011 2902 17075
rect 2966 17011 2967 17075
rect 2901 15416 2967 17011
rect 2901 15352 2902 15416
rect 2966 15352 2967 15416
rect 2901 13736 2967 15352
rect 2901 13672 2902 13736
rect 2966 13672 2967 13736
rect 2490 12742 2556 12743
rect 2490 12678 2491 12742
rect 2555 12678 2556 12742
rect 2490 12677 2556 12678
rect 696 11119 974 11183
rect 1038 11119 1044 11183
rect 696 1038 1044 11119
rect 2901 12056 2967 13672
rect 2901 11992 2902 12056
rect 2966 11992 2967 12056
rect 2901 10376 2967 11992
rect 2901 10312 2902 10376
rect 2966 10312 2967 10376
rect 2901 9468 2967 10312
rect 4005 21328 4071 22142
rect 4005 21264 4006 21328
rect 4070 21264 4071 21328
rect 4005 11183 4071 21264
rect 9630 19964 9706 22371
rect 10803 22353 10869 30787
rect 9630 19900 9636 19964
rect 9700 19900 9706 19964
rect 9630 19894 9706 19900
rect 10798 19815 10874 22353
rect 13305 20612 13381 20618
rect 13305 20548 13311 20612
rect 13375 20548 13381 20612
rect 12694 19822 12770 19828
rect 10798 19751 10804 19815
rect 10868 19751 10874 19815
rect 10798 19745 10874 19751
rect 12011 19815 12087 19821
rect 12011 19751 12017 19815
rect 12081 19751 12087 19815
rect 12011 19535 12087 19751
rect 12011 19471 12017 19535
rect 12081 19471 12087 19535
rect 12011 19465 12087 19471
rect 12694 19758 12700 19822
rect 12764 19758 12770 19822
rect 12694 19535 12770 19758
rect 12694 19471 12700 19535
rect 12764 19471 12770 19535
rect 12694 19465 12770 19471
rect 13305 19822 13381 20548
rect 13305 19758 13311 19822
rect 13375 19758 13381 19822
rect 13305 19535 13381 19758
rect 13305 19471 13311 19535
rect 13375 19471 13381 19535
rect 13305 18242 13381 19471
rect 13305 18178 13311 18242
rect 13375 18178 13381 18242
rect 13305 17452 13381 18178
rect 13730 20612 13806 20618
rect 13730 20548 13736 20612
rect 13800 20548 13806 20612
rect 13730 19822 13806 20548
rect 13730 19758 13736 19822
rect 13800 19758 13806 19822
rect 13730 18242 13806 19758
rect 14109 20605 14185 20611
rect 14109 20541 14115 20605
rect 14179 20541 14185 20605
rect 14109 19815 14185 20541
rect 14109 19751 14115 19815
rect 14179 19751 14185 19815
rect 14109 19535 14185 19751
rect 14109 19471 14115 19535
rect 14179 19471 14185 19535
rect 14109 19465 14185 19471
rect 16026 20419 16092 39989
rect 16026 20355 16027 20419
rect 16091 20355 16092 20419
rect 13730 18178 13736 18242
rect 13800 18178 13806 18242
rect 13730 18172 13806 18178
rect 14109 18235 14185 18241
rect 14109 18171 14115 18235
rect 14179 18171 14185 18235
rect 13305 17388 13311 17452
rect 13375 17388 13381 17452
rect 13305 15872 13381 17388
rect 13305 15808 13311 15872
rect 13375 15808 13381 15872
rect 13305 15082 13381 15808
rect 13730 17452 13806 17458
rect 13730 17388 13736 17452
rect 13800 17388 13806 17452
rect 13730 15872 13806 17388
rect 14109 17445 14185 18171
rect 14109 17381 14115 17445
rect 14179 17381 14185 17445
rect 14109 17375 14185 17381
rect 14505 18235 14581 18241
rect 14505 18171 14511 18235
rect 14575 18171 14581 18235
rect 14505 17445 14581 18171
rect 14505 17381 14511 17445
rect 14575 17381 14581 17445
rect 14505 17375 14581 17381
rect 13730 15808 13736 15872
rect 13800 15808 13806 15872
rect 13730 15802 13806 15808
rect 14109 15865 14185 15871
rect 5914 15075 5990 15081
rect 5914 15011 5920 15075
rect 5984 15011 5990 15075
rect 13305 15018 13311 15082
rect 13375 15018 13381 15082
rect 13305 15012 13381 15018
rect 14109 15801 14115 15865
rect 14179 15801 14185 15865
rect 14109 15075 14185 15801
rect 5914 12227 5990 15011
rect 14109 15011 14115 15075
rect 14179 15011 14185 15075
rect 14109 15005 14185 15011
rect 14505 15865 14581 15871
rect 14505 15801 14511 15865
rect 14575 15801 14581 15865
rect 14505 15075 14581 15801
rect 14505 15011 14511 15075
rect 14575 15011 14581 15075
rect 14505 15005 14581 15011
rect 16026 15027 16092 20355
rect 16026 14963 16027 15027
rect 16091 14963 16092 15027
rect 10714 14926 10790 14932
rect 10714 14862 10720 14926
rect 10784 14862 10790 14926
rect 10714 13641 10790 14862
rect 16026 14691 16092 14963
rect 16498 17445 16564 39989
rect 16498 17381 16499 17445
rect 16563 17381 16564 17445
rect 16498 14691 16564 17381
rect 4005 11119 4006 11183
rect 4070 11119 4071 11183
rect 4005 9612 4071 11119
rect 4005 9548 4006 9612
rect 4070 9548 4071 9612
rect 1570 8696 1646 8702
rect 1570 8632 1576 8696
rect 1640 8632 1646 8696
rect 1570 7016 1646 8632
rect 2896 8696 2972 9468
rect 4005 9409 4071 9548
rect 5919 9612 5985 12227
rect 5919 9548 5920 9612
rect 5984 9548 5985 9612
rect 2896 8632 2902 8696
rect 2966 8632 2972 8696
rect 2896 8626 2972 8632
rect 1570 6952 1576 7016
rect 1640 6952 1646 7016
rect 1570 5336 1646 6952
rect 1570 5272 1576 5336
rect 1640 5272 1646 5336
rect 1570 3656 1646 5272
rect 5919 3829 5985 9548
rect 10719 5243 10785 13641
rect 15440 12259 15516 12265
rect 15440 12195 15446 12259
rect 15510 12195 15516 12259
rect 15440 12046 15516 12195
rect 16021 12259 16097 14691
rect 16021 12195 16027 12259
rect 16091 12195 16097 12259
rect 16021 12189 16097 12195
rect 16493 14685 16569 14691
rect 16493 14621 16499 14685
rect 16563 14621 16569 14685
rect 16493 12073 16569 14621
rect 16930 14685 16996 39989
rect 16930 14621 16931 14685
rect 16995 14621 16996 14685
rect 16930 14615 16996 14621
rect 17274 15027 17340 39989
rect 17274 14963 17275 15027
rect 17339 14963 17340 15027
rect 17274 14615 17340 14963
rect 17698 14691 17764 39989
rect 18590 15027 18656 39991
rect 18590 14963 18591 15027
rect 18655 14963 18656 15027
rect 17693 14685 17769 14691
rect 17693 14621 17699 14685
rect 17763 14621 17769 14685
rect 17693 14489 17769 14621
rect 18590 14585 18656 14963
rect 19015 14659 19081 39993
rect 19658 15470 19724 39961
rect 19658 15406 19659 15470
rect 19723 15406 19724 15470
rect 19658 15027 19724 15406
rect 19658 14963 19659 15027
rect 19723 14963 19724 15027
rect 17693 14425 17699 14489
rect 17763 14425 17769 14489
rect 19010 14495 19086 14659
rect 19658 14615 19724 14963
rect 20906 14691 20972 39961
rect 19010 14431 19016 14495
rect 19080 14431 19086 14495
rect 19010 14425 19086 14431
rect 20901 14483 20977 14691
rect 17693 14419 17769 14425
rect 20901 14419 20907 14483
rect 20971 14419 20977 14483
rect 20901 14413 20977 14419
rect 22007 14483 22073 40642
rect 22007 14419 22008 14483
rect 22072 14419 22073 14483
rect 22007 13884 22073 14419
rect 22417 15470 22483 40642
rect 22417 15406 22418 15470
rect 22482 15406 22483 15470
rect 22417 13884 22483 15406
rect 45253 15055 45319 40642
rect 45253 14991 45254 15055
rect 45318 14991 45319 15055
rect 22002 13500 22078 13884
rect 21998 13494 22078 13500
rect 21998 13430 22004 13494
rect 22068 13430 22078 13494
rect 21998 13424 22078 13430
rect 15445 6378 15511 12046
rect 16493 11997 16726 12073
rect 6052 4338 6128 4344
rect 6052 4274 6058 4338
rect 6122 4274 6128 4338
rect 5733 3818 5990 3829
rect 5733 3754 5739 3818
rect 5803 3754 5990 3818
rect 5733 3753 5990 3754
rect 5733 3748 5809 3753
rect 1570 3592 1576 3656
rect 1640 3592 1646 3656
rect 1570 1976 1646 3592
rect 1570 1912 1576 1976
rect 1640 1912 1646 1976
rect 1570 1640 1646 1912
rect 1570 1576 1576 1640
rect 1640 1576 1646 1640
rect 1570 1570 1646 1576
rect 696 974 702 1038
rect 766 974 838 1038
rect 902 974 974 1038
rect 1038 974 1044 1038
rect 696 902 1044 974
rect 696 838 702 902
rect 766 838 838 902
rect 902 838 974 902
rect 1038 838 1044 902
rect 696 766 1044 838
rect 696 702 702 766
rect 766 702 838 766
rect 902 702 974 766
rect 1038 702 1044 766
rect 696 696 1044 702
rect 0 278 6 342
rect 70 278 142 342
rect 206 278 278 342
rect 342 278 348 342
rect 0 206 348 278
rect 0 142 6 206
rect 70 142 142 206
rect 206 142 278 206
rect 342 142 348 206
rect 0 70 348 142
rect 0 6 6 70
rect 70 6 142 70
rect 206 6 278 70
rect 342 6 348 70
rect 0 0 348 6
rect 6052 0 6128 4274
rect 10714 3894 10790 5243
rect 15440 4286 15516 6378
rect 16655 6351 16721 11997
rect 21998 11961 22074 11967
rect 21998 11897 22004 11961
rect 22068 11897 22074 11961
rect 21998 9745 22074 11897
rect 22412 11961 22488 13884
rect 45253 13808 45319 14991
rect 45663 40157 45729 40642
rect 45663 40093 45664 40157
rect 45728 40093 45729 40157
rect 45663 13808 45729 40093
rect 46759 40157 46835 40163
rect 46759 40093 46765 40157
rect 46829 40093 46835 40157
rect 49967 40151 50043 40157
rect 46759 39885 46835 40093
rect 48650 40145 48726 40151
rect 48650 40081 48656 40145
rect 48720 40081 48726 40145
rect 46764 14615 46830 39885
rect 48012 15055 48078 39961
rect 48650 39917 48726 40081
rect 49967 40087 49973 40151
rect 50037 40087 50043 40151
rect 48012 14991 48013 15055
rect 48077 14991 48078 15055
rect 48012 14615 48078 14991
rect 48655 14583 48721 39917
rect 49080 15055 49146 39991
rect 49967 39913 50043 40087
rect 49080 14991 49081 15055
rect 49145 14991 49146 15055
rect 49080 14585 49146 14991
rect 49972 14685 50038 39913
rect 49972 14621 49973 14685
rect 50037 14621 50038 14685
rect 49972 14615 50038 14621
rect 50396 15055 50462 39989
rect 50396 14991 50397 15055
rect 50461 14991 50462 15055
rect 50396 14615 50462 14991
rect 50740 14685 50806 39989
rect 51167 39913 51243 42453
rect 51639 42331 51715 42337
rect 51639 42267 51645 42331
rect 51709 42267 51715 42331
rect 51639 39913 51715 42267
rect 52220 42331 52296 42480
rect 52220 42267 52226 42331
rect 52290 42267 52296 42331
rect 52220 42261 52296 42267
rect 57035 42223 57101 47869
rect 61835 41012 61901 49283
rect 66174 49016 66250 50632
rect 66174 48952 66180 49016
rect 66244 48952 66250 49016
rect 63939 47944 64015 47950
rect 63939 47880 63945 47944
rect 64009 47880 64015 47944
rect 63939 47336 64015 47880
rect 63939 47272 63945 47336
rect 64009 47272 64015 47336
rect 63939 47266 64015 47272
rect 66174 47336 66250 48952
rect 66174 47272 66180 47336
rect 66244 47272 66250 47336
rect 66174 45656 66250 47272
rect 66174 45592 66180 45656
rect 66244 45592 66250 45656
rect 64848 43976 64924 43982
rect 64848 43912 64854 43976
rect 64918 43912 64924 43976
rect 61835 40948 61836 41012
rect 61900 40948 61901 41012
rect 61835 40809 61901 40948
rect 63749 41481 63815 43703
rect 64848 43644 64924 43912
rect 66174 43976 66250 45592
rect 66174 43912 66180 43976
rect 66244 43912 66250 43976
rect 66174 43906 66250 43912
rect 63749 41417 63750 41481
rect 63814 41417 63815 41481
rect 63749 41012 63815 41417
rect 63749 40948 63750 41012
rect 63814 40948 63815 41012
rect 50740 14621 50741 14685
rect 50805 14621 50806 14685
rect 50740 14615 50806 14621
rect 51172 18235 51238 39913
rect 51172 18171 51173 18235
rect 51237 18171 51238 18235
rect 51172 14685 51238 18171
rect 51172 14621 51173 14685
rect 51237 14621 51238 14685
rect 51172 14615 51238 14621
rect 51644 17259 51710 39913
rect 63749 31474 63815 40948
rect 63749 31410 63750 31474
rect 63814 31410 63815 31474
rect 63749 30970 63815 31410
rect 64853 42296 64919 43644
rect 64853 42232 64854 42296
rect 64918 42232 64919 42296
rect 64853 40616 64919 42232
rect 65264 41848 65330 41849
rect 65264 41784 65265 41848
rect 65329 41784 65330 41848
rect 65264 41783 65330 41784
rect 64853 40552 64854 40616
rect 64918 40552 64919 40616
rect 64853 38936 64919 40552
rect 64853 38872 64854 38936
rect 64918 38872 64919 38936
rect 64853 37163 64919 38872
rect 64853 37099 64854 37163
rect 64918 37099 64919 37163
rect 64853 35576 64919 37099
rect 64853 35512 64854 35576
rect 64918 35512 64919 35576
rect 64853 33896 64919 35512
rect 64853 33832 64854 33896
rect 64918 33832 64919 33896
rect 64853 32216 64919 33832
rect 64853 32152 64854 32216
rect 64918 32152 64919 32216
rect 64853 30987 64919 32152
rect 65267 31646 65327 41783
rect 66776 41481 67124 51700
rect 66776 41417 66782 41481
rect 66846 41417 67124 41481
rect 65264 31645 65330 31646
rect 65264 31581 65265 31645
rect 65329 31581 65330 31645
rect 65264 31580 65330 31581
rect 66776 31474 67124 41417
rect 66776 31410 66782 31474
rect 66846 31410 67124 31474
rect 63744 21328 63820 30970
rect 64848 30536 64924 30987
rect 64848 30472 64854 30536
rect 64918 30472 64924 30536
rect 64848 30466 64924 30472
rect 66174 30536 66250 30542
rect 66174 30472 66180 30536
rect 66244 30472 66250 30536
rect 66174 28856 66250 30472
rect 66174 28792 66180 28856
rect 66244 28792 66250 28856
rect 66174 27176 66250 28792
rect 66174 27112 66180 27176
rect 66244 27112 66250 27176
rect 66174 25496 66250 27112
rect 66174 25432 66180 25496
rect 66244 25432 66250 25496
rect 66174 23816 66250 25432
rect 66174 23752 66180 23816
rect 66244 23752 66250 23816
rect 66174 22136 66250 23752
rect 66174 22072 66180 22136
rect 66244 22072 66250 22136
rect 66174 22066 66250 22072
rect 63744 21264 63750 21328
rect 63814 21264 63820 21328
rect 63744 21258 63820 21264
rect 66776 21328 67124 31410
rect 66776 21264 66782 21328
rect 66846 21264 67124 21328
rect 54355 20612 54431 20618
rect 53155 20605 53231 20611
rect 53155 20541 53161 20605
rect 53225 20541 53231 20605
rect 53155 19815 53231 20541
rect 53155 19751 53161 19815
rect 53225 19751 53231 19815
rect 53155 19745 53231 19751
rect 53551 20605 53627 20611
rect 53551 20541 53557 20605
rect 53621 20541 53627 20605
rect 53551 19815 53627 20541
rect 54355 20548 54361 20612
rect 54425 20548 54431 20612
rect 53551 19751 53557 19815
rect 53621 19751 53627 19815
rect 53551 19535 53627 19751
rect 53551 19471 53557 19535
rect 53621 19471 53627 19535
rect 53551 18235 53627 19471
rect 53551 18171 53557 18235
rect 53621 18171 53627 18235
rect 53551 17732 53627 18171
rect 53551 17668 53557 17732
rect 53621 17668 53627 17732
rect 53551 17445 53627 17668
rect 53551 17381 53557 17445
rect 53621 17381 53627 17445
rect 53551 17375 53627 17381
rect 53930 19822 54006 19828
rect 53930 19758 53936 19822
rect 54000 19758 54006 19822
rect 53930 18242 54006 19758
rect 54355 19822 54431 20548
rect 54355 19758 54361 19822
rect 54425 19758 54431 19822
rect 54355 19535 54431 19758
rect 54355 19471 54361 19535
rect 54425 19471 54431 19535
rect 54355 19465 54431 19471
rect 66174 20456 66250 20462
rect 66174 20392 66180 20456
rect 66244 20392 66250 20456
rect 66174 18776 66250 20392
rect 66174 18712 66180 18776
rect 66244 18712 66250 18776
rect 53930 18178 53936 18242
rect 54000 18178 54006 18242
rect 53930 17452 54006 18178
rect 53930 17388 53936 17452
rect 54000 17388 54006 17452
rect 51644 17195 51645 17259
rect 51709 17195 51710 17259
rect 51644 15055 51710 17195
rect 53930 15872 54006 17388
rect 51644 14991 51645 15055
rect 51709 14991 51710 15055
rect 53155 15865 53231 15871
rect 53155 15801 53161 15865
rect 53225 15801 53231 15865
rect 53155 15075 53231 15801
rect 53155 15011 53161 15075
rect 53225 15011 53231 15075
rect 53155 15005 53231 15011
rect 53551 15865 53627 15871
rect 53551 15801 53557 15865
rect 53621 15801 53627 15865
rect 53930 15808 53936 15872
rect 54000 15808 54006 15872
rect 53930 15802 54006 15808
rect 54355 18242 54431 18248
rect 54355 18178 54361 18242
rect 54425 18178 54431 18242
rect 54355 17732 54431 18178
rect 54355 17668 54361 17732
rect 54425 17668 54431 17732
rect 54355 17452 54431 17668
rect 54355 17388 54361 17452
rect 54425 17388 54431 17452
rect 54355 15872 54431 17388
rect 54355 15808 54361 15872
rect 54425 15808 54431 15872
rect 53551 15075 53627 15801
rect 53551 15011 53557 15075
rect 53621 15011 53627 15075
rect 54355 15082 54431 15808
rect 54355 15018 54361 15082
rect 54425 15018 54431 15082
rect 66174 17096 66250 18712
rect 66174 17032 66180 17096
rect 66244 17032 66250 17096
rect 66174 15416 66250 17032
rect 66174 15352 66180 15416
rect 66244 15352 66250 15416
rect 54355 15012 54431 15018
rect 56946 15075 57022 15081
rect 53551 15005 53627 15011
rect 56946 15011 56952 15075
rect 57016 15011 57022 15075
rect 51644 14615 51710 14991
rect 56946 14623 57022 15011
rect 58114 14926 58190 14932
rect 58114 14862 58120 14926
rect 58184 14862 58190 14926
rect 22412 11897 22418 11961
rect 22482 11897 22488 11961
rect 22412 11891 22488 11897
rect 23628 13494 23704 13500
rect 23628 13430 23634 13494
rect 23698 13430 23704 13494
rect 21998 9681 22004 9745
rect 22068 9681 22074 9745
rect 21998 9675 22074 9681
rect 23490 9745 23566 9751
rect 23490 9681 23496 9745
rect 23560 9681 23566 9745
rect 21998 9308 22074 9314
rect 21998 9244 22004 9308
rect 22068 9244 22074 9308
rect 21998 8484 22074 9244
rect 23490 8976 23566 9681
rect 23628 9308 23704 13430
rect 23628 9244 23634 9308
rect 23698 9244 23704 9308
rect 23628 9238 23704 9244
rect 56951 11079 57017 14623
rect 58114 14605 58190 14862
rect 56951 11015 56952 11079
rect 57016 11015 57017 11079
rect 23490 8912 23496 8976
rect 23560 8912 23566 8976
rect 23490 8906 23566 8912
rect 40408 8976 40484 8982
rect 40408 8912 40414 8976
rect 40478 8912 40484 8976
rect 21998 8420 22004 8484
rect 22068 8420 22074 8484
rect 21998 8414 22074 8420
rect 15279 4210 15516 4286
rect 10714 3830 10720 3894
rect 10784 3830 10790 3894
rect 10714 3824 10790 3830
rect 11966 3894 12042 3900
rect 11966 3830 11972 3894
rect 12036 3830 12042 3894
rect 11966 1646 12042 3830
rect 14302 3894 14378 3900
rect 14302 3830 14308 3894
rect 14372 3830 14378 3894
rect 12136 3044 12212 3050
rect 12136 2980 12142 3044
rect 12206 2980 12212 3044
rect 11966 1640 12062 1646
rect 11966 1576 11992 1640
rect 12056 1576 12062 1640
rect 11966 1570 12062 1576
rect 12136 0 12212 2980
rect 13304 3044 13380 3050
rect 13304 2980 13310 3044
rect 13374 2980 13380 3044
rect 13134 2480 13210 2486
rect 13134 2416 13140 2480
rect 13204 2416 13210 2480
rect 13134 1038 13210 2416
rect 13134 974 13140 1038
rect 13204 974 13210 1038
rect 13134 968 13210 974
rect 13304 0 13380 2980
rect 14130 2480 14206 2486
rect 14130 2416 14136 2480
rect 14200 2416 14206 2480
rect 13666 1640 13742 1646
rect 13666 1576 13672 1640
rect 13736 1576 13742 1640
rect 13666 342 13742 1576
rect 14130 1038 14206 2416
rect 14302 1640 14378 3830
rect 14302 1576 14308 1640
rect 14372 1576 14378 1640
rect 14302 1570 14378 1576
rect 14472 3044 14548 3050
rect 14472 2980 14478 3044
rect 14542 2980 14548 3044
rect 14130 974 14136 1038
rect 14200 974 14206 1038
rect 14130 968 14206 974
rect 13666 278 13672 342
rect 13736 278 13742 342
rect 13666 272 13742 278
rect 14472 0 14548 2980
rect 15279 2480 15355 4210
rect 18706 3894 18782 3900
rect 18706 3830 18712 3894
rect 18776 3830 18782 3894
rect 15279 2416 15285 2480
rect 15349 2416 15355 2480
rect 15279 2410 15355 2416
rect 15640 3044 15716 3050
rect 15640 2980 15646 3044
rect 15710 2980 15716 3044
rect 15640 0 15716 2980
rect 16808 3044 16884 3050
rect 16808 2980 16814 3044
rect 16878 2980 16884 3044
rect 16808 0 16884 2980
rect 17976 3044 18052 3050
rect 17976 2980 17982 3044
rect 18046 2980 18052 3044
rect 17976 0 18052 2980
rect 18706 1640 18782 3830
rect 18706 1576 18712 1640
rect 18776 1576 18782 1640
rect 18706 1570 18782 1576
rect 19144 3044 19220 3050
rect 19144 2980 19150 3044
rect 19214 2980 19220 3044
rect 19144 0 19220 2980
rect 20312 3044 20388 3050
rect 20312 2980 20318 3044
rect 20382 2980 20388 3044
rect 20312 0 20388 2980
rect 21480 3044 21556 3050
rect 21480 2980 21486 3044
rect 21550 2980 21556 3044
rect 21480 0 21556 2980
rect 22648 3044 22724 3050
rect 22648 2980 22654 3044
rect 22718 2980 22724 3044
rect 22648 0 22724 2980
rect 27291 2480 27367 2486
rect 27291 2416 27297 2480
rect 27361 2416 27367 2480
rect 27106 1640 27182 1646
rect 27106 1576 27112 1640
rect 27176 1576 27182 1640
rect 27106 342 27182 1576
rect 27291 1038 27367 2416
rect 27291 974 27297 1038
rect 27361 974 27367 1038
rect 27291 968 27367 974
rect 40408 1038 40484 8912
rect 56951 6189 57017 11015
rect 57657 9588 57733 9594
rect 57657 9524 57663 9588
rect 57727 9524 57733 9588
rect 40408 974 40414 1038
rect 40478 974 40484 1038
rect 40408 968 40484 974
rect 40546 1640 40622 1646
rect 40546 1576 40552 1640
rect 40616 1576 40622 1640
rect 27106 278 27112 342
rect 27176 278 27182 342
rect 27106 272 27182 278
rect 40546 342 40622 1576
rect 40546 278 40552 342
rect 40616 278 40622 342
rect 40546 272 40622 278
rect 53986 1640 54062 1646
rect 53986 1576 53992 1640
rect 54056 1576 54062 1640
rect 53986 342 54062 1576
rect 56946 1038 57022 6189
rect 56946 974 56952 1038
rect 57016 974 57022 1038
rect 56946 968 57022 974
rect 53986 278 53992 342
rect 54056 278 54062 342
rect 53986 272 54062 278
rect 57657 0 57733 9524
rect 57795 8460 57871 8466
rect 57795 8396 57801 8460
rect 57865 8396 57871 8460
rect 57795 0 57871 8396
rect 57944 6760 58020 6766
rect 57944 6696 57950 6760
rect 58014 6696 58020 6760
rect 57944 0 58020 6696
rect 58119 6131 58185 14605
rect 66174 13736 66250 15352
rect 66174 13672 66180 13736
rect 66244 13672 66250 13736
rect 66174 12056 66250 13672
rect 66174 11992 66180 12056
rect 66244 11992 66250 12056
rect 66174 10376 66250 11992
rect 66174 10312 66180 10376
rect 66244 10312 66250 10376
rect 66174 8696 66250 10312
rect 66174 8632 66180 8696
rect 66244 8632 66250 8696
rect 66174 7016 66250 8632
rect 66174 6952 66180 7016
rect 66244 6952 66250 7016
rect 66174 5336 66250 6952
rect 66174 5272 66180 5336
rect 66244 5272 66250 5336
rect 66174 3656 66250 5272
rect 66174 3592 66180 3656
rect 66244 3592 66250 3656
rect 65746 1976 65822 1982
rect 65746 1912 65752 1976
rect 65816 1912 65822 1976
rect 65746 1640 65822 1912
rect 66174 1976 66250 3592
rect 66174 1912 66180 1976
rect 66244 1912 66250 1976
rect 66174 1906 66250 1912
rect 66776 11079 67124 21264
rect 66776 11015 66782 11079
rect 66846 11015 67124 11079
rect 65746 1576 65752 1640
rect 65816 1576 65822 1640
rect 65746 1570 65822 1576
rect 66776 1038 67124 11015
rect 66776 974 66782 1038
rect 66846 974 66918 1038
rect 66982 974 67054 1038
rect 67118 974 67124 1038
rect 66776 902 67124 974
rect 66776 838 66782 902
rect 66846 838 66918 902
rect 66982 838 67054 902
rect 67118 838 67124 902
rect 66776 766 67124 838
rect 66776 702 66782 766
rect 66846 702 66918 766
rect 66982 702 67054 766
rect 67118 702 67124 766
rect 66776 696 67124 702
rect 67472 42296 67820 52396
rect 67472 42232 67478 42296
rect 67542 42232 67820 42296
rect 67472 32216 67820 42232
rect 67472 32152 67478 32216
rect 67542 32152 67820 32216
rect 67472 22136 67820 32152
rect 67472 22072 67478 22136
rect 67542 22072 67820 22136
rect 67472 20456 67820 22072
rect 67472 20392 67478 20456
rect 67542 20392 67820 20456
rect 67472 10376 67820 20392
rect 67472 10312 67478 10376
rect 67542 10312 67820 10376
rect 67472 342 67820 10312
rect 67472 278 67478 342
rect 67542 278 67614 342
rect 67678 278 67750 342
rect 67814 278 67820 342
rect 67472 206 67820 278
rect 67472 142 67478 206
rect 67542 142 67614 206
rect 67678 142 67750 206
rect 67814 142 67820 206
rect 67472 70 67820 142
rect 67472 6 67478 70
rect 67542 6 67614 70
rect 67678 6 67750 70
rect 67814 6 67820 70
rect 67472 0 67820 6
use subbyte2_bank  subbyte2_bank_0
timestamp 1543373562
transform 1 0 11004 0 1 6302
box 0 0 45812 41924
use subbyte2_col_addr_dff  subbyte2_col_addr_dff_0
timestamp 1543373571
transform -1 0 54648 0 -1 50290
box -49 -49 2372 1467
use subbyte2_col_addr_dff  subbyte2_col_addr_dff_1
timestamp 1543373571
transform 1 0 12004 0 1 2448
box -49 -49 2372 1467
use subbyte2_contact_37  subbyte2_contact_37_0
timestamp 1543373572
transform 1 0 1512 0 1 51034
box 0 0 192 192
use subbyte2_contact_37  subbyte2_contact_37_1
timestamp 1543373572
transform 1 0 66116 0 1 51034
box 0 0 192 192
use subbyte2_contact_37  subbyte2_contact_37_2
timestamp 1543373572
transform 1 0 66116 0 1 1512
box 0 0 192 192
use subbyte2_contact_37  subbyte2_contact_37_3
timestamp 1543373572
transform 1 0 1512 0 1 1512
box 0 0 192 192
use subbyte2_control_logic_r  subbyte2_control_logic_r_0
timestamp 1543373571
transform -1 0 65254 0 -1 49326
box -75 -49 8270 18432
use subbyte2_control_logic_w  subbyte2_control_logic_w_0
timestamp 1543373571
transform 1 0 2566 0 1 3786
box -75 -49 8270 18432
use subbyte2_cr_3  subbyte2_cr_3_0
timestamp 1543373571
transform 1 0 11004 0 1 6302
box 2083 -3207 4411 2244
use subbyte2_cr_4  subbyte2_cr_4_0
timestamp 1543373571
transform 1 0 11004 0 1 6302
box 4376 -3230 30680 1874
use subbyte2_cr_5  subbyte2_cr_5_0
timestamp 1543373571
transform 1 0 11004 0 1 6302
box 41317 39678 42561 43341
use subbyte2_data_dff  subbyte2_data_dff_0
timestamp 1543373571
transform 1 0 14340 0 1 2448
box -49 -49 9380 1467
use subbyte2_row_addr_dff  subbyte2_row_addr_dff_0
timestamp 1543373571
transform -1 0 58152 0 -1 14648
box -75 -51 1243 8535
use subbyte2_row_addr_dff  subbyte2_row_addr_dff_1
timestamp 1543373571
transform 1 0 9668 0 1 22328
box -75 -51 1243 8535
<< labels >>
rlabel metal3 s 0 4312 76 4388 4 csb0
port 3 nsew
rlabel metal4 s 6052 0 6128 76 4 clk0
port 5 nsew
rlabel metal4 s 14472 0 14548 76 4 din0[0]
port 7 nsew
rlabel metal4 s 15640 0 15716 76 4 din0[1]
port 9 nsew
rlabel metal4 s 16808 0 16884 76 4 din0[2]
port 11 nsew
rlabel metal4 s 17976 0 18052 76 4 din0[3]
port 13 nsew
rlabel metal4 s 19144 0 19220 76 4 din0[4]
port 15 nsew
rlabel metal4 s 20312 0 20388 76 4 din0[5]
port 17 nsew
rlabel metal4 s 21480 0 21556 76 4 din0[6]
port 19 nsew
rlabel metal4 s 22648 0 22724 76 4 din0[7]
port 21 nsew
rlabel metal4 s 12136 0 12212 76 4 addr0[0]
port 23 nsew
rlabel metal4 s 13304 0 13380 76 4 addr0[1]
port 25 nsew
rlabel metal3 s 0 22854 76 22930 4 addr0[2]
port 27 nsew
rlabel metal3 s 0 24554 76 24630 4 addr0[3]
port 29 nsew
rlabel metal3 s 0 25682 76 25758 4 addr0[4]
port 31 nsew
rlabel metal3 s 0 27382 76 27458 4 addr0[5]
port 33 nsew
rlabel metal3 s 0 28510 76 28586 4 addr0[6]
port 35 nsew
rlabel metal3 s 0 30210 76 30286 4 addr0[7]
port 37 nsew
rlabel metal3 s 67744 48724 67820 48800 4 csb1
port 39 nsew
rlabel metal4 s 61692 52662 61768 52738 4 clk1
port 41 nsew
rlabel metal4 s 23973 52662 24049 52738 4 dout1[0]
port 43 nsew
rlabel metal4 s 26469 52662 26545 52738 4 dout1[1]
port 45 nsew
rlabel metal4 s 28965 52662 29041 52738 4 dout1[2]
port 47 nsew
rlabel metal4 s 31461 52662 31537 52738 4 dout1[3]
port 49 nsew
rlabel metal4 s 33957 52662 34033 52738 4 dout1[4]
port 51 nsew
rlabel metal4 s 36453 52662 36529 52738 4 dout1[5]
port 53 nsew
rlabel metal4 s 38949 52662 39025 52738 4 dout1[6]
port 55 nsew
rlabel metal4 s 41445 52662 41521 52738 4 dout1[7]
port 57 nsew
rlabel metal4 s 54440 52662 54516 52738 4 addr1[0]
port 59 nsew
rlabel metal4 s 53272 52662 53348 52738 4 addr1[1]
port 61 nsew
rlabel metal3 s 67744 14046 67820 14122 4 addr1[2]
port 63 nsew
rlabel metal3 s 67744 12346 67820 12422 4 addr1[3]
port 65 nsew
rlabel metal3 s 67744 11218 67820 11294 4 addr1[4]
port 67 nsew
rlabel metal4 s 57657 0 57733 76 4 addr1[5]
port 69 nsew
rlabel metal4 s 57795 0 57871 76 4 addr1[6]
port 71 nsew
rlabel metal4 s 57944 0 58020 76 4 addr1[7]
port 73 nsew
rlabel metal3 s 0 52390 67820 52738 4 vccd1
port 75 nsew
rlabel metal3 s 0 0 67820 348 4 vccd1
port 75 nsew
rlabel metal4 s 67472 0 67820 52738 4 vccd1
port 75 nsew
rlabel metal4 s 0 0 348 52738 4 vccd1
port 75 nsew
rlabel metal4 s 66776 696 67124 52042 4 vssd1
port 77 nsew
rlabel metal3 s 696 696 67124 1044 4 vssd1
port 77 nsew
rlabel metal3 s 696 51694 67124 52042 4 vssd1
port 77 nsew
rlabel metal4 s 696 696 1044 52042 4 vssd1
port 77 nsew
<< properties >>
string FIXED_BBOX 0 0 67820 52738
<< end >>
