magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1335 -1311 2503 9795
<< locali >>
rect 1151 8501 1185 8517
rect 1151 8451 1185 8467
rect -17 7087 17 7103
rect -17 7037 17 7053
rect 1151 5673 1185 5689
rect 1151 5623 1185 5639
rect -17 4259 17 4275
rect -17 4209 17 4225
rect 1151 2845 1185 2861
rect 1151 2795 1185 2811
rect -17 1431 17 1447
rect -17 1381 17 1397
rect 1151 17 1185 33
rect 1151 -33 1185 -17
<< viali >>
rect 1151 8467 1185 8501
rect -17 7053 17 7087
rect 1151 5639 1185 5673
rect -17 4225 17 4259
rect 1151 2811 1185 2845
rect -17 1397 17 1431
rect 1151 -17 1185 17
<< metal1 >>
rect 1136 8458 1142 8510
rect 1194 8458 1200 8510
rect -32 7044 -26 7096
rect 26 7044 32 7096
rect 1136 5630 1142 5682
rect 1194 5630 1200 5682
rect -32 4216 -26 4268
rect 26 4216 32 4268
rect 1136 2802 1142 2854
rect 1194 2802 1200 2854
rect -32 1388 -26 1440
rect 26 1388 32 1440
rect 1136 -26 1142 26
rect 1194 -26 1200 26
<< via1 >>
rect 1142 8501 1194 8510
rect 1142 8467 1151 8501
rect 1151 8467 1185 8501
rect 1185 8467 1194 8501
rect 1142 8458 1194 8467
rect -26 7087 26 7096
rect -26 7053 -17 7087
rect -17 7053 17 7087
rect 17 7053 26 7087
rect -26 7044 26 7053
rect 1142 5673 1194 5682
rect 1142 5639 1151 5673
rect 1151 5639 1185 5673
rect 1185 5639 1194 5673
rect 1142 5630 1194 5639
rect -26 4259 26 4268
rect -26 4225 -17 4259
rect -17 4225 17 4259
rect 17 4225 26 4259
rect -26 4216 26 4225
rect 1142 2845 1194 2854
rect 1142 2811 1151 2845
rect 1151 2811 1185 2845
rect 1185 2811 1194 2845
rect 1142 2802 1194 2811
rect -26 1431 26 1440
rect -26 1397 -17 1431
rect -17 1397 17 1431
rect 17 1397 26 1431
rect -26 1388 26 1397
rect 1142 17 1194 26
rect 1142 -17 1151 17
rect 1151 -17 1185 17
rect 1185 -17 1194 17
rect 1142 -26 1194 -17
<< metal2 >>
rect 1140 8512 1196 8521
rect 137 7894 203 7946
rect -28 7098 28 7107
rect -28 7033 28 7042
rect 137 6194 203 6246
rect 137 5066 203 5118
rect -28 4270 28 4279
rect -28 4205 28 4214
rect 137 3366 203 3418
rect 137 2238 203 2290
rect -28 1442 28 1451
rect -28 1377 28 1386
rect 137 538 203 590
rect 369 345 397 8484
rect 1140 8447 1196 8456
rect 1082 7823 1148 7875
rect 1082 6265 1148 6317
rect 1140 5684 1196 5693
rect 1140 5619 1196 5628
rect 1082 4995 1148 5047
rect 1082 3437 1148 3489
rect 1140 2856 1196 2865
rect 1140 2791 1196 2800
rect 1082 2167 1148 2219
rect 1082 609 1148 661
rect 368 336 424 345
rect 368 271 424 280
rect 369 0 397 271
rect 1140 28 1196 37
rect 1140 -37 1196 -28
<< via2 >>
rect 1140 8510 1196 8512
rect -28 7096 28 7098
rect -28 7044 -26 7096
rect -26 7044 26 7096
rect 26 7044 28 7096
rect -28 7042 28 7044
rect -28 4268 28 4270
rect -28 4216 -26 4268
rect -26 4216 26 4268
rect 26 4216 28 4268
rect -28 4214 28 4216
rect -28 1440 28 1442
rect -28 1388 -26 1440
rect -26 1388 26 1440
rect 26 1388 28 1440
rect -28 1386 28 1388
rect 1140 8458 1142 8510
rect 1142 8458 1194 8510
rect 1194 8458 1196 8510
rect 1140 8456 1196 8458
rect 1140 5682 1196 5684
rect 1140 5630 1142 5682
rect 1142 5630 1194 5682
rect 1194 5630 1196 5682
rect 1140 5628 1196 5630
rect 1140 2854 1196 2856
rect 1140 2802 1142 2854
rect 1142 2802 1194 2854
rect 1194 2802 1196 2854
rect 1140 2800 1196 2802
rect 368 280 424 336
rect 1140 26 1196 28
rect 1140 -26 1142 26
rect 1142 -26 1194 26
rect 1194 -26 1196 26
rect 1140 -28 1196 -26
<< metal3 >>
rect 1135 8516 1201 8517
rect 1093 8452 1136 8516
rect 1200 8452 1243 8516
rect 1135 8451 1201 8452
rect -33 7102 33 7103
rect -75 7038 -32 7102
rect 32 7038 75 7102
rect -33 7037 33 7038
rect 1135 5688 1201 5689
rect 1093 5624 1136 5688
rect 1200 5624 1243 5688
rect 1135 5623 1201 5624
rect -33 4274 33 4275
rect -75 4210 -32 4274
rect 32 4210 75 4274
rect -33 4209 33 4210
rect 1135 2860 1201 2861
rect 1093 2796 1136 2860
rect 1200 2796 1243 2860
rect 1135 2795 1201 2796
rect -33 1446 33 1447
rect -75 1382 -32 1446
rect 32 1382 75 1446
rect -33 1381 33 1382
rect 363 338 429 341
rect 0 336 1168 338
rect 0 280 368 336
rect 424 280 1168 336
rect 0 278 1168 280
rect 363 275 429 278
rect 1135 32 1201 33
rect 1093 -32 1136 32
rect 1200 -32 1243 32
rect 1135 -33 1201 -32
<< via3 >>
rect 1136 8512 1200 8516
rect 1136 8456 1140 8512
rect 1140 8456 1196 8512
rect 1196 8456 1200 8512
rect 1136 8452 1200 8456
rect -32 7098 32 7102
rect -32 7042 -28 7098
rect -28 7042 28 7098
rect 28 7042 32 7098
rect -32 7038 32 7042
rect 1136 5684 1200 5688
rect 1136 5628 1140 5684
rect 1140 5628 1196 5684
rect 1196 5628 1200 5684
rect 1136 5624 1200 5628
rect -32 4270 32 4274
rect -32 4214 -28 4270
rect -28 4214 28 4270
rect 28 4214 32 4270
rect -32 4210 32 4214
rect 1136 2856 1200 2860
rect 1136 2800 1140 2856
rect 1140 2800 1196 2856
rect 1196 2800 1200 2856
rect 1136 2796 1200 2800
rect -32 1442 32 1446
rect -32 1386 -28 1442
rect -28 1386 28 1442
rect 28 1386 32 1442
rect -32 1382 32 1386
rect 1136 28 1200 32
rect 1136 -28 1140 28
rect 1140 -28 1196 28
rect 1196 -28 1200 28
rect 1136 -32 1200 -28
<< metal4 >>
rect -33 7102 33 8517
rect -33 7038 -32 7102
rect 32 7038 33 7102
rect -33 4274 33 7038
rect -33 4210 -32 4274
rect 32 4210 33 4274
rect -33 1446 33 4210
rect -33 1382 -32 1446
rect 32 1382 33 1446
rect -33 -33 33 1382
rect 1135 8516 1201 8535
rect 1135 8452 1136 8516
rect 1200 8452 1201 8516
rect 1135 5688 1201 8452
rect 1135 5624 1136 5688
rect 1200 5624 1201 5688
rect 1135 2860 1201 5624
rect 1135 2796 1136 2860
rect 1200 2796 1201 2860
rect 1135 32 1201 2796
rect 1135 -32 1136 32
rect 1200 -32 1201 32
rect 1135 -51 1201 -32
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1438349329
transform 1 0 0 0 -1 8484
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1438349329
transform 1 0 0 0 1 5656
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1438349329
transform 1 0 0 0 -1 5656
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1438349329
transform 1 0 0 0 1 2828
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_4
timestamp 1438349329
transform 1 0 0 0 -1 2828
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_5
timestamp 1438349329
transform 1 0 0 0 1 0
box -36 -43 1204 1467
<< labels >>
rlabel metal4 s -33 -33 33 8517 4 vdd
port 3 nsew
rlabel metal4 s 1135 -51 1201 8535 4 gnd
port 5 nsew
rlabel metal2 s 137 538 203 590 4 din_0
port 7 nsew
rlabel metal2 s 1082 609 1148 661 4 dout_0
port 9 nsew
rlabel metal2 s 137 2238 203 2290 4 din_1
port 11 nsew
rlabel metal2 s 1082 2167 1148 2219 4 dout_1
port 13 nsew
rlabel metal2 s 137 3366 203 3418 4 din_2
port 15 nsew
rlabel metal2 s 1082 3437 1148 3489 4 dout_2
port 17 nsew
rlabel metal2 s 137 5066 203 5118 4 din_3
port 19 nsew
rlabel metal2 s 1082 4995 1148 5047 4 dout_3
port 21 nsew
rlabel metal2 s 137 6194 203 6246 4 din_4
port 23 nsew
rlabel metal2 s 1082 6265 1148 6317 4 dout_4
port 25 nsew
rlabel metal2 s 137 7894 203 7946 4 din_5
port 27 nsew
rlabel metal2 s 1082 7823 1148 7875 4 dout_5
port 29 nsew
rlabel metal3 s 0 278 1168 338 4 clk
port 31 nsew
<< properties >>
string FIXED_BBOX 1135 -37 1201 -33
<< end >>
