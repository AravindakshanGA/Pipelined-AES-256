magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect 3116 -4490 31940 3134
<< metal1 >>
rect 13101 1811 13107 1863
rect 13159 1811 13165 1863
rect 15597 1811 15603 1863
rect 15655 1811 15661 1863
rect 18093 1811 18099 1863
rect 18151 1811 18157 1863
rect 20589 1811 20595 1863
rect 20647 1811 20653 1863
rect 23085 1811 23091 1863
rect 23143 1811 23149 1863
rect 25581 1811 25587 1863
rect 25639 1811 25645 1863
rect 28077 1811 28083 1863
rect 28135 1811 28141 1863
rect 30573 1811 30579 1863
rect 30631 1811 30637 1863
<< via1 >>
rect 13107 1811 13159 1863
rect 15603 1811 15655 1863
rect 18099 1811 18151 1863
rect 20595 1811 20647 1863
rect 23091 1811 23143 1863
rect 25587 1811 25639 1863
rect 28083 1811 28135 1863
rect 30579 1811 30631 1863
<< metal2 >>
rect 13105 1865 13161 1874
rect 13105 1800 13161 1809
rect 15601 1865 15657 1874
rect 15601 1800 15657 1809
rect 18097 1865 18153 1874
rect 18097 1800 18153 1809
rect 20593 1865 20649 1874
rect 20593 1800 20649 1809
rect 23089 1865 23145 1874
rect 23089 1800 23145 1809
rect 25585 1865 25641 1874
rect 25585 1800 25641 1809
rect 28081 1865 28137 1874
rect 28081 1800 28137 1809
rect 30577 1865 30633 1874
rect 30577 1800 30633 1809
rect 4423 -3165 4479 -3156
rect 4423 -3230 4479 -3221
rect 5591 -3165 5647 -3156
rect 5591 -3230 5647 -3221
rect 6759 -3165 6815 -3156
rect 6759 -3230 6815 -3221
rect 7927 -3165 7983 -3156
rect 7927 -3230 7983 -3221
rect 9095 -3165 9151 -3156
rect 9095 -3230 9151 -3221
rect 10263 -3165 10319 -3156
rect 10263 -3230 10319 -3221
rect 11431 -3165 11487 -3156
rect 11431 -3230 11487 -3221
rect 12599 -3165 12655 -3156
rect 12599 -3230 12655 -3221
<< via2 >>
rect 13105 1863 13161 1865
rect 13105 1811 13107 1863
rect 13107 1811 13159 1863
rect 13159 1811 13161 1863
rect 13105 1809 13161 1811
rect 15601 1863 15657 1865
rect 15601 1811 15603 1863
rect 15603 1811 15655 1863
rect 15655 1811 15657 1863
rect 15601 1809 15657 1811
rect 18097 1863 18153 1865
rect 18097 1811 18099 1863
rect 18099 1811 18151 1863
rect 18151 1811 18153 1863
rect 18097 1809 18153 1811
rect 20593 1863 20649 1865
rect 20593 1811 20595 1863
rect 20595 1811 20647 1863
rect 20647 1811 20649 1863
rect 20593 1809 20649 1811
rect 23089 1863 23145 1865
rect 23089 1811 23091 1863
rect 23091 1811 23143 1863
rect 23143 1811 23145 1863
rect 23089 1809 23145 1811
rect 25585 1863 25641 1865
rect 25585 1811 25587 1863
rect 25587 1811 25639 1863
rect 25639 1811 25641 1863
rect 25585 1809 25641 1811
rect 28081 1863 28137 1865
rect 28081 1811 28083 1863
rect 28083 1811 28135 1863
rect 28135 1811 28137 1863
rect 28081 1809 28137 1811
rect 30577 1863 30633 1865
rect 30577 1811 30579 1863
rect 30579 1811 30631 1863
rect 30631 1811 30633 1863
rect 30577 1809 30633 1811
rect 4423 -3221 4479 -3165
rect 5591 -3221 5647 -3165
rect 6759 -3221 6815 -3165
rect 7927 -3221 7983 -3165
rect 9095 -3221 9151 -3165
rect 10263 -3221 10319 -3165
rect 11431 -3221 11487 -3165
rect 12599 -3221 12655 -3165
<< metal3 >>
rect 13100 1869 13166 1870
rect 15596 1869 15662 1870
rect 18092 1869 18158 1870
rect 20588 1869 20654 1870
rect 23084 1869 23150 1870
rect 25580 1869 25646 1870
rect 28076 1869 28142 1870
rect 30572 1869 30638 1870
rect 13058 1805 13101 1869
rect 13165 1805 13208 1869
rect 15554 1805 15597 1869
rect 15661 1805 15704 1869
rect 18050 1805 18093 1869
rect 18157 1805 18200 1869
rect 20546 1805 20589 1869
rect 20653 1805 20696 1869
rect 23042 1805 23085 1869
rect 23149 1805 23192 1869
rect 25538 1805 25581 1869
rect 25645 1805 25688 1869
rect 28034 1805 28077 1869
rect 28141 1805 28184 1869
rect 30530 1805 30573 1869
rect 30637 1805 30680 1869
rect 13100 1804 13166 1805
rect 15596 1804 15662 1805
rect 18092 1804 18158 1805
rect 20588 1804 20654 1805
rect 23084 1804 23150 1805
rect 25580 1804 25646 1805
rect 28076 1804 28142 1805
rect 30572 1804 30638 1805
rect 12589 -516 12595 -452
rect 12659 -454 12665 -452
rect 30567 -454 30573 -452
rect 12659 -514 30573 -454
rect 12659 -516 12665 -514
rect 30567 -516 30573 -514
rect 30637 -516 30643 -452
rect 11421 -760 11427 -696
rect 11491 -698 11497 -696
rect 28071 -698 28077 -696
rect 11491 -758 28077 -698
rect 11491 -760 11497 -758
rect 28071 -760 28077 -758
rect 28141 -760 28147 -696
rect 10253 -1004 10259 -940
rect 10323 -942 10329 -940
rect 25575 -942 25581 -940
rect 10323 -1002 25581 -942
rect 10323 -1004 10329 -1002
rect 25575 -1004 25581 -1002
rect 25645 -1004 25651 -940
rect 9085 -1248 9091 -1184
rect 9155 -1186 9161 -1184
rect 23079 -1186 23085 -1184
rect 9155 -1246 23085 -1186
rect 9155 -1248 9161 -1246
rect 23079 -1248 23085 -1246
rect 23149 -1248 23155 -1184
rect 7917 -1492 7923 -1428
rect 7987 -1430 7993 -1428
rect 20583 -1430 20589 -1428
rect 7987 -1490 20589 -1430
rect 7987 -1492 7993 -1490
rect 20583 -1492 20589 -1490
rect 20653 -1492 20659 -1428
rect 6749 -1736 6755 -1672
rect 6819 -1674 6825 -1672
rect 18087 -1674 18093 -1672
rect 6819 -1734 18093 -1674
rect 6819 -1736 6825 -1734
rect 18087 -1736 18093 -1734
rect 18157 -1736 18163 -1672
rect 5581 -1980 5587 -1916
rect 5651 -1918 5657 -1916
rect 15591 -1918 15597 -1916
rect 5651 -1978 15597 -1918
rect 5651 -1980 5657 -1978
rect 15591 -1980 15597 -1978
rect 15661 -1980 15667 -1916
rect 4413 -2224 4419 -2160
rect 4483 -2162 4489 -2160
rect 13095 -2162 13101 -2160
rect 4483 -2222 13101 -2162
rect 4483 -2224 4489 -2222
rect 13095 -2224 13101 -2222
rect 13165 -2224 13171 -2160
rect 4418 -3161 4484 -3160
rect 5586 -3161 5652 -3160
rect 6754 -3161 6820 -3160
rect 7922 -3161 7988 -3160
rect 9090 -3161 9156 -3160
rect 10258 -3161 10324 -3160
rect 11426 -3161 11492 -3160
rect 12594 -3161 12660 -3160
rect 4376 -3225 4419 -3161
rect 4483 -3225 4526 -3161
rect 5544 -3225 5587 -3161
rect 5651 -3225 5694 -3161
rect 6712 -3225 6755 -3161
rect 6819 -3225 6862 -3161
rect 7880 -3225 7923 -3161
rect 7987 -3225 8030 -3161
rect 9048 -3225 9091 -3161
rect 9155 -3225 9198 -3161
rect 10216 -3225 10259 -3161
rect 10323 -3225 10366 -3161
rect 11384 -3225 11427 -3161
rect 11491 -3225 11534 -3161
rect 12552 -3225 12595 -3161
rect 12659 -3225 12702 -3161
rect 4418 -3226 4484 -3225
rect 5586 -3226 5652 -3225
rect 6754 -3226 6820 -3225
rect 7922 -3226 7988 -3225
rect 9090 -3226 9156 -3225
rect 10258 -3226 10324 -3225
rect 11426 -3226 11492 -3225
rect 12594 -3226 12660 -3225
<< via3 >>
rect 13101 1865 13165 1869
rect 13101 1809 13105 1865
rect 13105 1809 13161 1865
rect 13161 1809 13165 1865
rect 13101 1805 13165 1809
rect 15597 1865 15661 1869
rect 15597 1809 15601 1865
rect 15601 1809 15657 1865
rect 15657 1809 15661 1865
rect 15597 1805 15661 1809
rect 18093 1865 18157 1869
rect 18093 1809 18097 1865
rect 18097 1809 18153 1865
rect 18153 1809 18157 1865
rect 18093 1805 18157 1809
rect 20589 1865 20653 1869
rect 20589 1809 20593 1865
rect 20593 1809 20649 1865
rect 20649 1809 20653 1865
rect 20589 1805 20653 1809
rect 23085 1865 23149 1869
rect 23085 1809 23089 1865
rect 23089 1809 23145 1865
rect 23145 1809 23149 1865
rect 23085 1805 23149 1809
rect 25581 1865 25645 1869
rect 25581 1809 25585 1865
rect 25585 1809 25641 1865
rect 25641 1809 25645 1865
rect 25581 1805 25645 1809
rect 28077 1865 28141 1869
rect 28077 1809 28081 1865
rect 28081 1809 28137 1865
rect 28137 1809 28141 1865
rect 28077 1805 28141 1809
rect 30573 1865 30637 1869
rect 30573 1809 30577 1865
rect 30577 1809 30633 1865
rect 30633 1809 30637 1865
rect 30573 1805 30637 1809
rect 12595 -516 12659 -452
rect 30573 -516 30637 -452
rect 11427 -760 11491 -696
rect 28077 -760 28141 -696
rect 10259 -1004 10323 -940
rect 25581 -1004 25645 -940
rect 9091 -1248 9155 -1184
rect 23085 -1248 23149 -1184
rect 7923 -1492 7987 -1428
rect 20589 -1492 20653 -1428
rect 6755 -1736 6819 -1672
rect 18093 -1736 18157 -1672
rect 5587 -1980 5651 -1916
rect 15597 -1980 15661 -1916
rect 4419 -2224 4483 -2160
rect 13101 -2224 13165 -2160
rect 4419 -3165 4483 -3161
rect 4419 -3221 4423 -3165
rect 4423 -3221 4479 -3165
rect 4479 -3221 4483 -3165
rect 4419 -3225 4483 -3221
rect 5587 -3165 5651 -3161
rect 5587 -3221 5591 -3165
rect 5591 -3221 5647 -3165
rect 5647 -3221 5651 -3165
rect 5587 -3225 5651 -3221
rect 6755 -3165 6819 -3161
rect 6755 -3221 6759 -3165
rect 6759 -3221 6815 -3165
rect 6815 -3221 6819 -3165
rect 6755 -3225 6819 -3221
rect 7923 -3165 7987 -3161
rect 7923 -3221 7927 -3165
rect 7927 -3221 7983 -3165
rect 7983 -3221 7987 -3165
rect 7923 -3225 7987 -3221
rect 9091 -3165 9155 -3161
rect 9091 -3221 9095 -3165
rect 9095 -3221 9151 -3165
rect 9151 -3221 9155 -3165
rect 9091 -3225 9155 -3221
rect 10259 -3165 10323 -3161
rect 10259 -3221 10263 -3165
rect 10263 -3221 10319 -3165
rect 10319 -3221 10323 -3165
rect 10259 -3225 10323 -3221
rect 11427 -3165 11491 -3161
rect 11427 -3221 11431 -3165
rect 11431 -3221 11487 -3165
rect 11487 -3221 11491 -3165
rect 11427 -3225 11491 -3221
rect 12595 -3165 12659 -3161
rect 12595 -3221 12599 -3165
rect 12599 -3221 12655 -3165
rect 12655 -3221 12659 -3165
rect 12595 -3225 12659 -3221
<< metal4 >>
rect 13100 1869 13166 1870
rect 13100 1805 13101 1869
rect 13165 1805 13166 1869
rect 13100 1804 13166 1805
rect 15596 1869 15662 1870
rect 15596 1805 15597 1869
rect 15661 1805 15662 1869
rect 15596 1804 15662 1805
rect 18092 1869 18158 1870
rect 18092 1805 18093 1869
rect 18157 1805 18158 1869
rect 18092 1804 18158 1805
rect 20588 1869 20654 1870
rect 20588 1805 20589 1869
rect 20653 1805 20654 1869
rect 20588 1804 20654 1805
rect 23084 1869 23150 1870
rect 23084 1805 23085 1869
rect 23149 1805 23150 1869
rect 23084 1804 23150 1805
rect 25580 1869 25646 1870
rect 25580 1805 25581 1869
rect 25645 1805 25646 1869
rect 25580 1804 25646 1805
rect 28076 1869 28142 1870
rect 28076 1805 28077 1869
rect 28141 1805 28142 1869
rect 28076 1804 28142 1805
rect 30572 1869 30638 1870
rect 30572 1805 30573 1869
rect 30637 1805 30638 1869
rect 30572 1804 30638 1805
rect 12594 -452 12660 -451
rect 12594 -516 12595 -452
rect 12659 -516 12660 -452
rect 12594 -517 12660 -516
rect 11426 -696 11492 -695
rect 11426 -760 11427 -696
rect 11491 -760 11492 -696
rect 11426 -761 11492 -760
rect 10258 -940 10324 -939
rect 10258 -1004 10259 -940
rect 10323 -1004 10324 -940
rect 10258 -1005 10324 -1004
rect 9090 -1184 9156 -1183
rect 9090 -1248 9091 -1184
rect 9155 -1248 9156 -1184
rect 9090 -1249 9156 -1248
rect 7922 -1428 7988 -1427
rect 7922 -1492 7923 -1428
rect 7987 -1492 7988 -1428
rect 7922 -1493 7988 -1492
rect 6754 -1672 6820 -1671
rect 6754 -1736 6755 -1672
rect 6819 -1736 6820 -1672
rect 6754 -1737 6820 -1736
rect 5586 -1916 5652 -1915
rect 5586 -1980 5587 -1916
rect 5651 -1980 5652 -1916
rect 5586 -1981 5652 -1980
rect 4418 -2160 4484 -2159
rect 4418 -2224 4419 -2160
rect 4483 -2224 4484 -2160
rect 4418 -2225 4484 -2224
rect 4421 -3160 4481 -2225
rect 5589 -3160 5649 -1981
rect 6757 -3160 6817 -1737
rect 7925 -3160 7985 -1493
rect 9093 -3160 9153 -1249
rect 10261 -3160 10321 -1005
rect 11429 -3160 11489 -761
rect 12597 -3160 12657 -517
rect 13103 -2159 13163 1804
rect 15599 -1915 15659 1804
rect 18095 -1671 18155 1804
rect 20591 -1427 20651 1804
rect 23087 -1183 23147 1804
rect 25583 -939 25643 1804
rect 28079 -695 28139 1804
rect 30575 -451 30635 1804
rect 30572 -452 30638 -451
rect 30572 -516 30573 -452
rect 30637 -516 30638 -452
rect 30572 -517 30638 -516
rect 28076 -696 28142 -695
rect 28076 -760 28077 -696
rect 28141 -760 28142 -696
rect 28076 -761 28142 -760
rect 25580 -940 25646 -939
rect 25580 -1004 25581 -940
rect 25645 -1004 25646 -940
rect 25580 -1005 25646 -1004
rect 23084 -1184 23150 -1183
rect 23084 -1248 23085 -1184
rect 23149 -1248 23150 -1184
rect 23084 -1249 23150 -1248
rect 20588 -1428 20654 -1427
rect 20588 -1492 20589 -1428
rect 20653 -1492 20654 -1428
rect 20588 -1493 20654 -1492
rect 18092 -1672 18158 -1671
rect 18092 -1736 18093 -1672
rect 18157 -1736 18158 -1672
rect 18092 -1737 18158 -1736
rect 15596 -1916 15662 -1915
rect 15596 -1980 15597 -1916
rect 15661 -1980 15662 -1916
rect 15596 -1981 15662 -1980
rect 13100 -2160 13166 -2159
rect 13100 -2224 13101 -2160
rect 13165 -2224 13166 -2160
rect 13100 -2225 13166 -2224
rect 4418 -3161 4484 -3160
rect 4418 -3225 4419 -3161
rect 4483 -3225 4484 -3161
rect 4418 -3226 4484 -3225
rect 5586 -3161 5652 -3160
rect 5586 -3225 5587 -3161
rect 5651 -3225 5652 -3161
rect 5586 -3226 5652 -3225
rect 6754 -3161 6820 -3160
rect 6754 -3225 6755 -3161
rect 6819 -3225 6820 -3161
rect 6754 -3226 6820 -3225
rect 7922 -3161 7988 -3160
rect 7922 -3225 7923 -3161
rect 7987 -3225 7988 -3161
rect 7922 -3226 7988 -3225
rect 9090 -3161 9156 -3160
rect 9090 -3225 9091 -3161
rect 9155 -3225 9156 -3161
rect 9090 -3226 9156 -3225
rect 10258 -3161 10324 -3160
rect 10258 -3225 10259 -3161
rect 10323 -3225 10324 -3161
rect 10258 -3226 10324 -3225
rect 11426 -3161 11492 -3160
rect 11426 -3225 11427 -3161
rect 11491 -3225 11492 -3161
rect 11426 -3226 11492 -3225
rect 12594 -3161 12660 -3160
rect 12594 -3225 12595 -3161
rect 12659 -3225 12660 -3161
rect 12594 -3226 12660 -3225
<< properties >>
string FIXED_BBOX 4376 -3230 30680 1874
<< end >>
