magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1335 -1309 9530 19692
<< locali >>
rect 8169 9915 8203 9931
rect 5634 9881 8169 9915
rect 8169 9865 8203 9881
rect 4801 9208 4835 9224
rect 3450 9171 3484 9187
rect 4801 9158 4835 9174
rect 3450 9121 3484 9137
rect 3369 8501 3403 8517
rect 3403 8467 5634 8501
rect 3369 8451 3403 8467
rect 3450 7832 3484 7848
rect 3450 7782 3484 7798
rect 3565 7832 3599 7848
rect 3565 7782 3599 7798
rect 8169 7087 8203 7103
rect 3754 7053 8169 7087
rect 8169 7037 8203 7053
rect 3733 6790 3952 6824
rect 3918 6308 3952 6790
rect 5573 6380 5607 6396
rect 5573 6330 5607 6346
rect 3598 6191 3632 6207
rect 3598 6141 3632 6157
rect 3498 5943 3532 5959
rect 3498 5893 3532 5909
rect 3369 5673 3403 5689
rect 3403 5639 6082 5673
rect 3369 5623 3403 5639
rect 3465 5403 3499 5419
rect 3465 5353 3499 5369
rect 3598 5279 3632 5295
rect 3598 5229 3632 5245
rect 3731 5155 3765 5171
rect 3731 5105 3765 5121
rect 4477 4966 4511 4982
rect 4477 4916 4511 4932
rect 8169 4259 8203 4275
rect 4780 4225 8169 4259
rect 8169 4209 8203 4225
rect 4269 3536 4303 3552
rect 4269 3486 4303 3502
rect 3598 3363 3632 3379
rect 3598 3313 3632 3329
rect 3498 3115 3532 3131
rect 3498 3065 3532 3081
rect 3369 2845 3403 2861
rect 3403 2811 5148 2845
rect 3369 2795 3403 2811
rect 3715 2541 3900 2575
rect 3450 2176 3484 2192
rect 3715 2176 3749 2541
rect 3966 2327 4000 2343
rect 3966 2277 4000 2293
rect 3582 2142 3749 2176
rect 4637 2154 4671 2170
rect 3450 2126 3484 2142
rect 4637 2104 4671 2120
rect 8169 1431 8203 1447
rect 5148 1397 8169 1431
rect 8169 1381 8203 1397
rect 7029 724 7063 740
rect 3450 686 3484 702
rect 7029 674 7063 690
rect 3450 636 3484 652
rect 3369 17 3403 33
rect 3403 -17 8186 17
rect 3369 -33 3403 -17
<< viali >>
rect 8169 9881 8203 9915
rect 3450 9137 3484 9171
rect 4801 9174 4835 9208
rect 3369 8467 3403 8501
rect 3450 7798 3484 7832
rect 3565 7798 3599 7832
rect 8169 7053 8203 7087
rect 5573 6346 5607 6380
rect 3598 6157 3632 6191
rect 3498 5909 3532 5943
rect 3369 5639 3403 5673
rect 3465 5369 3499 5403
rect 3598 5245 3632 5279
rect 3731 5121 3765 5155
rect 4477 4932 4511 4966
rect 8169 4225 8203 4259
rect 4269 3502 4303 3536
rect 3598 3329 3632 3363
rect 3498 3081 3532 3115
rect 3369 2811 3403 2845
rect 3966 2293 4000 2327
rect 3450 2142 3484 2176
rect 4637 2120 4671 2154
rect 8169 1397 8203 1431
rect 3450 652 3484 686
rect 7029 690 7063 724
rect 3369 -17 3403 17
<< metal1 >>
rect 8154 9872 8160 9924
rect 8212 9872 8218 9924
rect 2948 9128 2954 9180
rect 3006 9168 3012 9180
rect 3438 9171 3496 9177
rect 3438 9168 3450 9171
rect 3006 9140 3450 9168
rect 3006 9128 3012 9140
rect 3438 9137 3450 9140
rect 3484 9137 3496 9171
rect 4786 9165 4792 9217
rect 4844 9165 4850 9217
rect 3438 9131 3496 9137
rect 3354 8458 3360 8510
rect 3412 8458 3418 8510
rect 2864 7789 2870 7841
rect 2922 7829 2928 7841
rect 3438 7832 3496 7838
rect 3438 7829 3450 7832
rect 2922 7801 3450 7829
rect 2922 7789 2928 7801
rect 3438 7798 3450 7801
rect 3484 7798 3496 7832
rect 3438 7792 3496 7798
rect 3550 7789 3556 7841
rect 3608 7789 3614 7841
rect 8154 7044 8160 7096
rect 8212 7044 8218 7096
rect 5558 6337 5564 6389
rect 5616 6337 5622 6389
rect 2864 6148 2870 6200
rect 2922 6188 2928 6200
rect 3586 6191 3644 6197
rect 3586 6188 3598 6191
rect 2922 6160 3598 6188
rect 2922 6148 2928 6160
rect 3586 6157 3598 6160
rect 3632 6157 3644 6191
rect 3586 6151 3644 6157
rect 3032 5900 3038 5952
rect 3090 5940 3096 5952
rect 3486 5943 3544 5949
rect 3486 5940 3498 5943
rect 3090 5912 3498 5940
rect 3090 5900 3096 5912
rect 3486 5909 3498 5912
rect 3532 5909 3544 5943
rect 3486 5903 3544 5909
rect 3354 5630 3360 5682
rect 3412 5630 3418 5682
rect 3200 5360 3206 5412
rect 3258 5400 3264 5412
rect 3453 5403 3511 5409
rect 3453 5400 3465 5403
rect 3258 5372 3465 5400
rect 3258 5360 3264 5372
rect 3453 5369 3465 5372
rect 3499 5369 3511 5403
rect 3453 5363 3511 5369
rect 2780 5236 2786 5288
rect 2838 5276 2844 5288
rect 3586 5279 3644 5285
rect 3586 5276 3598 5279
rect 2838 5248 3598 5276
rect 2838 5236 2844 5248
rect 3586 5245 3598 5248
rect 3632 5245 3644 5279
rect 3586 5239 3644 5245
rect 2948 5112 2954 5164
rect 3006 5152 3012 5164
rect 3719 5155 3777 5161
rect 3719 5152 3731 5155
rect 3006 5124 3731 5152
rect 3006 5112 3012 5124
rect 3719 5121 3731 5124
rect 3765 5121 3777 5155
rect 3719 5115 3777 5121
rect 4462 4923 4468 4975
rect 4520 4923 4526 4975
rect 1521 4296 1527 4348
rect 1579 4336 1585 4348
rect 2864 4336 2870 4348
rect 1579 4308 2870 4336
rect 1579 4296 1585 4308
rect 2864 4296 2870 4308
rect 2922 4296 2928 4348
rect 8154 4216 8160 4268
rect 8212 4216 8218 4268
rect 351 4136 357 4188
rect 409 4176 415 4188
rect 3116 4176 3122 4188
rect 409 4148 3122 4176
rect 409 4136 415 4148
rect 3116 4136 3122 4148
rect 3174 4136 3180 4188
rect 4254 3493 4260 3545
rect 4312 3493 4318 3545
rect 3200 3320 3206 3372
rect 3258 3360 3264 3372
rect 3586 3363 3644 3369
rect 3586 3360 3598 3363
rect 3258 3332 3598 3360
rect 3258 3320 3264 3332
rect 3586 3329 3598 3332
rect 3632 3329 3644 3363
rect 3586 3323 3644 3329
rect 3116 3072 3122 3124
rect 3174 3112 3180 3124
rect 3486 3115 3544 3121
rect 3486 3112 3498 3115
rect 3174 3084 3498 3112
rect 3174 3072 3180 3084
rect 3486 3081 3498 3084
rect 3532 3081 3544 3115
rect 3486 3075 3544 3081
rect 3354 2802 3360 2854
rect 3412 2802 3418 2854
rect 3951 2284 3957 2336
rect 4009 2284 4015 2336
rect 3116 2133 3122 2185
rect 3174 2173 3180 2185
rect 3438 2176 3496 2182
rect 3438 2173 3450 2176
rect 3174 2145 3450 2173
rect 3174 2133 3180 2145
rect 3438 2142 3450 2145
rect 3484 2142 3496 2176
rect 3438 2136 3496 2142
rect 4622 2111 4628 2163
rect 4680 2111 4686 2163
rect 8154 1388 8160 1440
rect 8212 1388 8218 1440
rect 3435 643 3441 695
rect 3493 643 3499 695
rect 7014 681 7020 733
rect 7072 681 7078 733
rect 3354 -26 3360 26
rect 3412 -26 3418 26
<< via1 >>
rect 8160 9915 8212 9924
rect 8160 9881 8169 9915
rect 8169 9881 8203 9915
rect 8203 9881 8212 9915
rect 8160 9872 8212 9881
rect 2954 9128 3006 9180
rect 4792 9208 4844 9217
rect 4792 9174 4801 9208
rect 4801 9174 4835 9208
rect 4835 9174 4844 9208
rect 4792 9165 4844 9174
rect 3360 8501 3412 8510
rect 3360 8467 3369 8501
rect 3369 8467 3403 8501
rect 3403 8467 3412 8501
rect 3360 8458 3412 8467
rect 2870 7789 2922 7841
rect 3556 7832 3608 7841
rect 3556 7798 3565 7832
rect 3565 7798 3599 7832
rect 3599 7798 3608 7832
rect 3556 7789 3608 7798
rect 8160 7087 8212 7096
rect 8160 7053 8169 7087
rect 8169 7053 8203 7087
rect 8203 7053 8212 7087
rect 8160 7044 8212 7053
rect 5564 6380 5616 6389
rect 5564 6346 5573 6380
rect 5573 6346 5607 6380
rect 5607 6346 5616 6380
rect 5564 6337 5616 6346
rect 2870 6148 2922 6200
rect 3038 5900 3090 5952
rect 3360 5673 3412 5682
rect 3360 5639 3369 5673
rect 3369 5639 3403 5673
rect 3403 5639 3412 5673
rect 3360 5630 3412 5639
rect 3206 5360 3258 5412
rect 2786 5236 2838 5288
rect 2954 5112 3006 5164
rect 4468 4966 4520 4975
rect 4468 4932 4477 4966
rect 4477 4932 4511 4966
rect 4511 4932 4520 4966
rect 4468 4923 4520 4932
rect 1527 4296 1579 4348
rect 2870 4296 2922 4348
rect 8160 4259 8212 4268
rect 8160 4225 8169 4259
rect 8169 4225 8203 4259
rect 8203 4225 8212 4259
rect 8160 4216 8212 4225
rect 357 4136 409 4188
rect 3122 4136 3174 4188
rect 4260 3536 4312 3545
rect 4260 3502 4269 3536
rect 4269 3502 4303 3536
rect 4303 3502 4312 3536
rect 4260 3493 4312 3502
rect 3206 3320 3258 3372
rect 3122 3072 3174 3124
rect 3360 2845 3412 2854
rect 3360 2811 3369 2845
rect 3369 2811 3403 2845
rect 3403 2811 3412 2845
rect 3360 2802 3412 2811
rect 3957 2327 4009 2336
rect 3957 2293 3966 2327
rect 3966 2293 4000 2327
rect 4000 2293 4009 2327
rect 3957 2284 4009 2293
rect 3122 2133 3174 2185
rect 4628 2154 4680 2163
rect 4628 2120 4637 2154
rect 4637 2120 4671 2154
rect 4671 2120 4680 2154
rect 4628 2111 4680 2120
rect 8160 1431 8212 1440
rect 8160 1397 8169 1431
rect 8169 1397 8203 1431
rect 8203 1397 8212 1431
rect 8160 1388 8212 1397
rect 3441 686 3493 695
rect 3441 652 3450 686
rect 3450 652 3484 686
rect 3484 652 3493 686
rect 3441 643 3493 652
rect 7020 724 7072 733
rect 7020 690 7029 724
rect 7029 690 7063 724
rect 7063 690 7072 724
rect 7020 681 7072 690
rect 3360 17 3412 26
rect 3360 -17 3369 17
rect 3369 -17 3403 17
rect 3403 -17 3412 17
rect 3360 -26 3412 -17
<< metal2 >>
rect -57 17699 -29 17727
rect 2798 7428 2826 9938
rect 2882 7847 2910 9938
rect 2966 9186 2994 9938
rect 2954 9180 3006 9186
rect 2954 9122 3006 9128
rect 2870 7841 2922 7847
rect 2870 7783 2922 7789
rect 2784 7419 2840 7428
rect 2784 7354 2840 7363
rect 1539 4354 1567 6401
rect 2798 5294 2826 7354
rect 2882 6206 2910 7783
rect 2870 6200 2922 6206
rect 2870 6142 2922 6148
rect 2786 5288 2838 5294
rect 2786 5230 2838 5236
rect 1527 4348 1579 4354
rect 1527 4290 1579 4296
rect 357 4188 409 4194
rect 357 4130 409 4136
rect 369 1414 397 4130
rect 1844 913 1900 922
rect 1844 848 1900 857
rect 137 538 203 590
rect 2798 0 2826 5230
rect 2882 4354 2910 6142
rect 2966 5170 2994 9122
rect 3050 5958 3078 9938
rect 3038 5952 3090 5958
rect 3038 5894 3090 5900
rect 2954 5164 3006 5170
rect 2954 5106 3006 5112
rect 2870 4348 2922 4354
rect 2870 4290 2922 4296
rect 2882 0 2910 4290
rect 2966 1750 2994 5106
rect 3050 3556 3078 5894
rect 3134 4194 3162 9938
rect 3218 5418 3246 9938
rect 8158 9926 8214 9935
rect 8158 9861 8214 9870
rect 4792 9217 4844 9223
rect 4844 9177 8270 9205
rect 4792 9159 4844 9165
rect 3358 8512 3414 8521
rect 3358 8447 3414 8456
rect 3556 7841 3608 7847
rect 3556 7783 3608 7789
rect 3568 7428 3596 7783
rect 3554 7419 3610 7428
rect 3554 7354 3610 7363
rect 8158 7098 8214 7107
rect 8158 7033 8214 7042
rect 5564 6389 5616 6395
rect 5616 6349 8270 6377
rect 5564 6331 5616 6337
rect 3358 5684 3414 5693
rect 3358 5619 3414 5628
rect 3206 5412 3258 5418
rect 3206 5354 3258 5360
rect 3122 4188 3174 4194
rect 3122 4130 3174 4136
rect 3036 3547 3092 3556
rect 3036 3482 3092 3491
rect 2952 1741 3008 1750
rect 2952 1676 3008 1685
rect 2966 0 2994 1676
rect 3050 0 3078 3482
rect 3134 3130 3162 4130
rect 3218 3378 3246 5354
rect 4468 4975 4520 4981
rect 4520 4935 8270 4963
rect 4468 4917 4520 4923
rect 8158 4270 8214 4279
rect 8158 4205 8214 4214
rect 4258 3547 4314 3556
rect 4258 3482 4314 3491
rect 3206 3372 3258 3378
rect 3206 3314 3258 3320
rect 3122 3124 3174 3130
rect 3122 3066 3174 3072
rect 3134 2191 3162 3066
rect 3218 2347 3246 3314
rect 3358 2856 3414 2865
rect 3358 2791 3414 2800
rect 3204 2338 3260 2347
rect 3204 2273 3260 2282
rect 3955 2338 4011 2347
rect 3955 2273 4011 2282
rect 3122 2185 3174 2191
rect 3122 2127 3174 2133
rect 3134 320 3162 2127
rect 3218 922 3246 2273
rect 4628 2163 4680 2169
rect 4628 2105 4680 2111
rect 4640 1750 4668 2105
rect 4626 1741 4682 1750
rect 4626 1676 4682 1685
rect 8158 1442 8214 1451
rect 8158 1377 8214 1386
rect 3204 913 3260 922
rect 3204 848 3260 857
rect 3120 311 3176 320
rect 3120 246 3176 255
rect 3134 0 3162 246
rect 3218 0 3246 848
rect 7020 733 7072 739
rect 3441 695 3493 701
rect 7072 693 8270 721
rect 7020 675 7072 681
rect 3441 637 3493 643
rect 7032 320 7060 675
rect 7018 311 7074 320
rect 7018 246 7074 255
rect 3358 28 3414 37
rect 3358 -37 3414 -28
<< via2 >>
rect 2784 7363 2840 7419
rect 1844 857 1900 913
rect 8158 9924 8214 9926
rect 8158 9872 8160 9924
rect 8160 9872 8212 9924
rect 8212 9872 8214 9924
rect 8158 9870 8214 9872
rect 3358 8510 3414 8512
rect 3358 8458 3360 8510
rect 3360 8458 3412 8510
rect 3412 8458 3414 8510
rect 3358 8456 3414 8458
rect 3554 7363 3610 7419
rect 8158 7096 8214 7098
rect 8158 7044 8160 7096
rect 8160 7044 8212 7096
rect 8212 7044 8214 7096
rect 8158 7042 8214 7044
rect 3358 5682 3414 5684
rect 3358 5630 3360 5682
rect 3360 5630 3412 5682
rect 3412 5630 3414 5682
rect 3358 5628 3414 5630
rect 3036 3491 3092 3547
rect 2952 1685 3008 1741
rect 8158 4268 8214 4270
rect 8158 4216 8160 4268
rect 8160 4216 8212 4268
rect 8212 4216 8214 4268
rect 8158 4214 8214 4216
rect 4258 3545 4314 3547
rect 4258 3493 4260 3545
rect 4260 3493 4312 3545
rect 4312 3493 4314 3545
rect 4258 3491 4314 3493
rect 3358 2854 3414 2856
rect 3358 2802 3360 2854
rect 3360 2802 3412 2854
rect 3412 2802 3414 2854
rect 3358 2800 3414 2802
rect 3204 2282 3260 2338
rect 3955 2336 4011 2338
rect 3955 2284 3957 2336
rect 3957 2284 4009 2336
rect 4009 2284 4011 2336
rect 3955 2282 4011 2284
rect 4626 1685 4682 1741
rect 8158 1440 8214 1442
rect 8158 1388 8160 1440
rect 8160 1388 8212 1440
rect 8212 1388 8214 1440
rect 8158 1386 8214 1388
rect 3204 857 3260 913
rect 3120 255 3176 311
rect 7018 255 7074 311
rect 3358 26 3414 28
rect 3358 -26 3360 26
rect 3360 -26 3412 26
rect 3412 -26 3414 26
rect 3358 -28 3414 -26
<< metal3 >>
rect 8153 9930 8219 9931
rect 8111 9866 8154 9930
rect 8218 9866 8261 9930
rect 8153 9865 8219 9866
rect 3353 8516 3419 8517
rect 3311 8452 3354 8516
rect 3418 8452 3461 8516
rect 3353 8451 3419 8452
rect 2779 7421 2845 7424
rect 3549 7421 3615 7424
rect 2779 7419 3615 7421
rect 2779 7363 2784 7419
rect 2840 7363 3554 7419
rect 3610 7363 3615 7419
rect 2779 7361 3615 7363
rect 2779 7358 2845 7361
rect 3549 7358 3615 7361
rect 8153 7102 8219 7103
rect 8111 7038 8154 7102
rect 8218 7038 8261 7102
rect 8153 7037 8219 7038
rect 3353 5688 3419 5689
rect 3311 5624 3354 5688
rect 3418 5624 3461 5688
rect 3353 5623 3419 5624
rect 8153 4274 8219 4275
rect 8111 4210 8154 4274
rect 8218 4210 8261 4274
rect 8153 4209 8219 4210
rect 3031 3549 3097 3552
rect 4253 3549 4319 3552
rect 3031 3547 4319 3549
rect 3031 3491 3036 3547
rect 3092 3491 4258 3547
rect 4314 3491 4319 3547
rect 3031 3489 4319 3491
rect 3031 3486 3097 3489
rect 4253 3486 4319 3489
rect 3353 2860 3419 2861
rect 3311 2796 3354 2860
rect 3418 2796 3461 2860
rect 3353 2795 3419 2796
rect 3199 2340 3265 2343
rect 3950 2340 4016 2343
rect 3199 2338 4016 2340
rect 3199 2282 3204 2338
rect 3260 2282 3955 2338
rect 4011 2282 4016 2338
rect 3199 2280 4016 2282
rect 3199 2277 3265 2280
rect 3950 2277 4016 2280
rect 2947 1743 3013 1746
rect 4621 1743 4687 1746
rect 2947 1741 4687 1743
rect 2947 1685 2952 1741
rect 3008 1685 4626 1741
rect 4682 1685 4687 1741
rect 2947 1683 4687 1685
rect 2947 1680 3013 1683
rect 4621 1680 4687 1683
rect 1228 1365 1326 1463
rect 8153 1446 8219 1447
rect 8111 1382 8154 1446
rect 8218 1382 8261 1446
rect 8153 1381 8219 1382
rect 1839 915 1905 918
rect 3199 915 3265 918
rect 1839 913 3265 915
rect 1839 857 1844 913
rect 1900 857 3204 913
rect 3260 857 3265 913
rect 1839 855 3265 857
rect 1839 852 1905 855
rect 3199 852 3265 855
rect 3115 313 3181 316
rect 7013 313 7079 316
rect 3115 311 7079 313
rect 3115 255 3120 311
rect 3176 255 7018 311
rect 7074 255 7079 311
rect 3115 253 7079 255
rect 3115 250 3181 253
rect 7013 250 7079 253
rect 1228 -49 1326 49
rect 3353 32 3419 33
rect 3311 -32 3354 32
rect 3418 -32 3461 32
rect 3353 -33 3419 -32
<< via3 >>
rect 8154 9926 8218 9930
rect 8154 9870 8158 9926
rect 8158 9870 8214 9926
rect 8214 9870 8218 9926
rect 8154 9866 8218 9870
rect 3354 8512 3418 8516
rect 3354 8456 3358 8512
rect 3358 8456 3414 8512
rect 3414 8456 3418 8512
rect 3354 8452 3418 8456
rect 8154 7098 8218 7102
rect 8154 7042 8158 7098
rect 8158 7042 8214 7098
rect 8214 7042 8218 7098
rect 8154 7038 8218 7042
rect 3354 5684 3418 5688
rect 3354 5628 3358 5684
rect 3358 5628 3414 5684
rect 3414 5628 3418 5684
rect 3354 5624 3418 5628
rect 8154 4270 8218 4274
rect 8154 4214 8158 4270
rect 8158 4214 8214 4270
rect 8214 4214 8218 4270
rect 8154 4210 8218 4214
rect 3354 2856 3418 2860
rect 3354 2800 3358 2856
rect 3358 2800 3414 2856
rect 3414 2800 3418 2856
rect 3354 2796 3418 2800
rect 8154 1442 8218 1446
rect 8154 1386 8158 1442
rect 8158 1386 8214 1442
rect 8214 1386 8218 1442
rect 8154 1382 8218 1386
rect 3354 28 3418 32
rect 3354 -28 3358 28
rect 3358 -28 3414 28
rect 3414 -28 3418 28
rect 3354 -32 3418 -28
<< metal4 >>
rect 335 5606 401 18415
rect 1439 5623 1505 18432
rect 8153 9930 8219 9931
rect 8153 9866 8154 9930
rect 8218 9866 8219 9930
rect 3353 8516 3419 8517
rect 3353 8452 3354 8516
rect 3418 8452 3419 8516
rect 3353 5688 3419 8452
rect 3353 5624 3354 5688
rect 3418 5624 3419 5688
rect 3353 2860 3419 5624
rect 3353 2796 3354 2860
rect 3418 2796 3419 2860
rect 3353 32 3419 2796
rect 8153 7102 8219 9866
rect 8153 7038 8154 7102
rect 8218 7038 8219 7102
rect 8153 4274 8219 7038
rect 8153 4210 8154 4274
rect 8218 4210 8219 4274
rect 8153 1446 8219 4210
rect 8153 1382 8154 1446
rect 8218 1382 8219 1446
rect 8153 1381 8219 1382
rect 3353 -32 3354 32
rect 3418 -32 3419 32
rect 3353 -33 3419 -32
use subbyte2_delay_chain  subbyte2_delay_chain_0
timestamp 1543373571
transform 1 0 0 0 -1 18382
box -75 -50 1876 12783
use subbyte2_dff_buf_array  subbyte2_dff_buf_array_0
timestamp 1543373571
transform 1 0 0 0 1 0
box -36 -49 2590 1471
use subbyte2_pand2_0  subbyte2_pand2_0_0
timestamp 1543373571
transform 1 0 3386 0 1 2828
box -36 -17 1430 1471
use subbyte2_pand2_0  subbyte2_pand2_0_1
timestamp 1543373571
transform 1 0 3754 0 -1 2828
box -36 -17 1430 1471
use subbyte2_pand3  subbyte2_pand3_0
timestamp 1543373571
transform 1 0 3386 0 -1 5656
box -36 -17 1746 1471
use subbyte2_pdriver_1  subbyte2_pdriver_1_0
timestamp 1543373571
transform 1 0 3386 0 1 0
box -36 -17 4836 1471
use subbyte2_pdriver_2  subbyte2_pdriver_2_0
timestamp 1543373571
transform 1 0 3386 0 1 8484
box -36 -17 2284 1471
use subbyte2_pdriver_5  subbyte2_pdriver_5_0
timestamp 1543373571
transform 1 0 3854 0 1 5656
box -36 -17 2264 1471
use subbyte2_pinv_0  subbyte2_pinv_0_0
timestamp 1543373571
transform 1 0 3386 0 -1 8484
box -36 -17 404 1471
use subbyte2_pinv_0  subbyte2_pinv_0_1
timestamp 1543373571
transform 1 0 3386 0 -1 2828
box -36 -17 404 1471
use subbyte2_pnand2_0  subbyte2_pnand2_0_0
timestamp 1543373571
transform 1 0 3386 0 1 5656
box -36 -17 504 1471
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
port 3 nsew
rlabel metal2 s 4818 9177 8270 9205 4 wl_en
port 5 nsew
rlabel metal2 s 4494 4935 8270 4963 4 w_en
port 7 nsew
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
port 9 nsew
rlabel metal2 s 5590 6349 8270 6377 4 p_en_bar
port 11 nsew
rlabel metal2 s 3453 655 3481 683 4 clk
port 13 nsew
rlabel metal2 s 7046 693 8270 721 4 clk_buf
port 15 nsew
rlabel metal4 s 335 5606 401 18415 4 vdd
port 17 nsew
rlabel metal3 s 1228 1365 1326 1463 4 vdd
port 17 nsew
rlabel metal4 s 8153 1381 8219 9931 4 vdd
port 17 nsew
rlabel metal4 s 3353 -33 3419 8517 4 gnd
port 19 nsew
rlabel metal3 s 1228 -49 1326 49 4 gnd
port 19 nsew
rlabel metal4 s 1439 5623 1505 18432 4 gnd
port 19 nsew
<< properties >>
string FIXED_BBOX 3353 -37 3419 -33
<< end >>
