magic
tech sky130A
magscale 1 2
timestamp 1543373569
<< checkpaint >>
rect -1260 -841 1926 27701
<< metal2 >>
rect 330 26015 438 26125
rect 0 25919 28 25967
rect 330 25795 438 25871
rect 0 25699 28 25747
rect 0 25603 28 25651
rect 330 25479 438 25555
rect 0 25383 28 25431
rect 330 25225 438 25335
rect 0 25129 28 25177
rect 330 25005 438 25081
rect 0 24909 28 24957
rect 0 24813 28 24861
rect 330 24689 438 24765
rect 0 24593 28 24641
rect 330 24435 438 24545
rect 0 24339 28 24387
rect 330 24215 438 24291
rect 0 24119 28 24167
rect 0 24023 28 24071
rect 330 23899 438 23975
rect 0 23803 28 23851
rect 330 23645 438 23755
rect 0 23549 28 23597
rect 330 23425 438 23501
rect 0 23329 28 23377
rect 0 23233 28 23281
rect 330 23109 438 23185
rect 0 23013 28 23061
rect 330 22855 438 22965
rect 0 22759 28 22807
rect 330 22635 438 22711
rect 0 22539 28 22587
rect 0 22443 28 22491
rect 330 22319 438 22395
rect 0 22223 28 22271
rect 330 22065 438 22175
rect 0 21969 28 22017
rect 330 21845 438 21921
rect 0 21749 28 21797
rect 0 21653 28 21701
rect 330 21529 438 21605
rect 0 21433 28 21481
rect 330 21275 438 21385
rect 0 21179 28 21227
rect 330 21055 438 21131
rect 0 20959 28 21007
rect 0 20863 28 20911
rect 330 20739 438 20815
rect 0 20643 28 20691
rect 330 20485 438 20595
rect 0 20389 28 20437
rect 330 20265 438 20341
rect 0 20169 28 20217
rect 0 20073 28 20121
rect 330 19949 438 20025
rect 0 19853 28 19901
rect 330 19695 438 19805
rect 0 19599 28 19647
rect 330 19475 438 19551
rect 0 19379 28 19427
rect 0 19283 28 19331
rect 330 19159 438 19235
rect 0 19063 28 19111
rect 330 18905 438 19015
rect 0 18809 28 18857
rect 330 18685 438 18761
rect 0 18589 28 18637
rect 0 18493 28 18541
rect 330 18369 438 18445
rect 0 18273 28 18321
rect 330 18115 438 18225
rect 0 18019 28 18067
rect 330 17895 438 17971
rect 0 17799 28 17847
rect 0 17703 28 17751
rect 330 17579 438 17655
rect 0 17483 28 17531
rect 330 17325 438 17435
rect 0 17229 28 17277
rect 330 17105 438 17181
rect 0 17009 28 17057
rect 0 16913 28 16961
rect 330 16789 438 16865
rect 0 16693 28 16741
rect 330 16535 438 16645
rect 0 16439 28 16487
rect 330 16315 438 16391
rect 0 16219 28 16267
rect 0 16123 28 16171
rect 330 15999 438 16075
rect 0 15903 28 15951
rect 330 15745 438 15855
rect 0 15649 28 15697
rect 330 15525 438 15601
rect 0 15429 28 15477
rect 0 15333 28 15381
rect 330 15209 438 15285
rect 0 15113 28 15161
rect 330 14955 438 15065
rect 0 14859 28 14907
rect 330 14735 438 14811
rect 0 14639 28 14687
rect 0 14543 28 14591
rect 330 14419 438 14495
rect 0 14323 28 14371
rect 330 14165 438 14275
rect 0 14069 28 14117
rect 330 13945 438 14021
rect 0 13849 28 13897
rect 0 13753 28 13801
rect 330 13629 438 13705
rect 0 13533 28 13581
rect 330 13375 438 13485
rect 0 13279 28 13327
rect 330 13155 438 13231
rect 0 13059 28 13107
rect 0 12963 28 13011
rect 330 12839 438 12915
rect 0 12743 28 12791
rect 330 12585 438 12695
rect 0 12489 28 12537
rect 330 12365 438 12441
rect 0 12269 28 12317
rect 0 12173 28 12221
rect 330 12049 438 12125
rect 0 11953 28 12001
rect 330 11795 438 11905
rect 0 11699 28 11747
rect 330 11575 438 11651
rect 0 11479 28 11527
rect 0 11383 28 11431
rect 330 11259 438 11335
rect 0 11163 28 11211
rect 330 11005 438 11115
rect 0 10909 28 10957
rect 330 10785 438 10861
rect 0 10689 28 10737
rect 0 10593 28 10641
rect 330 10469 438 10545
rect 0 10373 28 10421
rect 330 10215 438 10325
rect 0 10119 28 10167
rect 330 9995 438 10071
rect 0 9899 28 9947
rect 0 9803 28 9851
rect 330 9679 438 9755
rect 0 9583 28 9631
rect 330 9425 438 9535
rect 0 9329 28 9377
rect 330 9205 438 9281
rect 0 9109 28 9157
rect 0 9013 28 9061
rect 330 8889 438 8965
rect 0 8793 28 8841
rect 330 8635 438 8745
rect 0 8539 28 8587
rect 330 8415 438 8491
rect 0 8319 28 8367
rect 0 8223 28 8271
rect 330 8099 438 8175
rect 0 8003 28 8051
rect 330 7845 438 7955
rect 0 7749 28 7797
rect 330 7625 438 7701
rect 0 7529 28 7577
rect 0 7433 28 7481
rect 330 7309 438 7385
rect 0 7213 28 7261
rect 330 7055 438 7165
rect 0 6959 28 7007
rect 330 6835 438 6911
rect 0 6739 28 6787
rect 0 6643 28 6691
rect 330 6519 438 6595
rect 0 6423 28 6471
rect 330 6265 438 6375
rect 0 6169 28 6217
rect 330 6045 438 6121
rect 0 5949 28 5997
rect 0 5853 28 5901
rect 330 5729 438 5805
rect 0 5633 28 5681
rect 330 5475 438 5585
rect 0 5379 28 5427
rect 330 5255 438 5331
rect 0 5159 28 5207
rect 0 5063 28 5111
rect 330 4939 438 5015
rect 0 4843 28 4891
rect 330 4685 438 4795
rect 0 4589 28 4637
rect 330 4465 438 4541
rect 0 4369 28 4417
rect 0 4273 28 4321
rect 330 4149 438 4225
rect 0 4053 28 4101
rect 330 3895 438 4005
rect 0 3799 28 3847
rect 330 3675 438 3751
rect 0 3579 28 3627
rect 0 3483 28 3531
rect 330 3359 438 3435
rect 0 3263 28 3311
rect 330 3105 438 3215
rect 0 3009 28 3057
rect 330 2885 438 2961
rect 0 2789 28 2837
rect 0 2693 28 2741
rect 330 2569 438 2645
rect 0 2473 28 2521
rect 330 2315 438 2425
rect 0 2219 28 2267
rect 330 2095 438 2171
rect 0 1999 28 2047
rect 0 1903 28 1951
rect 330 1779 438 1855
rect 0 1683 28 1731
rect 330 1525 438 1635
rect 0 1429 28 1477
rect 330 1305 438 1381
rect 0 1209 28 1257
rect 0 1113 28 1161
rect 330 989 438 1065
rect 0 893 28 941
rect 330 735 438 845
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_0
timestamp -19799
transform -1 0 624 0 1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_1
timestamp -19799
transform -1 0 624 0 -1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_2
timestamp -19799
transform -1 0 624 0 1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_3
timestamp -19799
transform -1 0 624 0 -1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_4
timestamp -19799
transform -1 0 624 0 1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_5
timestamp -19799
transform -1 0 624 0 -1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_6
timestamp -19799
transform -1 0 624 0 1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_7
timestamp -19799
transform -1 0 624 0 -1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_8
timestamp -19799
transform -1 0 624 0 1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_9
timestamp -19799
transform -1 0 624 0 -1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_10
timestamp -19799
transform -1 0 624 0 1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_11
timestamp -19799
transform -1 0 624 0 -1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_12
timestamp -19799
transform -1 0 624 0 1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_13
timestamp -19799
transform -1 0 624 0 -1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_14
timestamp -19799
transform -1 0 624 0 1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_15
timestamp -19799
transform -1 0 624 0 -1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_16
timestamp -19799
transform -1 0 624 0 1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_17
timestamp -19799
transform -1 0 624 0 -1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_18
timestamp -19799
transform -1 0 624 0 1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_19
timestamp -19799
transform -1 0 624 0 -1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_20
timestamp -19799
transform -1 0 624 0 1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_21
timestamp -19799
transform -1 0 624 0 -1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_22
timestamp -19799
transform -1 0 624 0 1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_23
timestamp -19799
transform -1 0 624 0 -1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_24
timestamp -19799
transform -1 0 624 0 1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_25
timestamp -19799
transform -1 0 624 0 -1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_26
timestamp -19799
transform -1 0 624 0 1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_27
timestamp -19799
transform -1 0 624 0 -1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_28
timestamp -19799
transform -1 0 624 0 1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_29
timestamp -19799
transform -1 0 624 0 -1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_30
timestamp -19799
transform -1 0 624 0 1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_31
timestamp -19799
transform -1 0 624 0 -1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_32
timestamp -19799
transform -1 0 624 0 1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_33
timestamp -19799
transform -1 0 624 0 -1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_34
timestamp -19799
transform -1 0 624 0 1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_35
timestamp -19799
transform -1 0 624 0 -1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_36
timestamp -19799
transform -1 0 624 0 1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_37
timestamp -19799
transform -1 0 624 0 -1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_38
timestamp -19799
transform -1 0 624 0 1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_39
timestamp -19799
transform -1 0 624 0 -1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_40
timestamp -19799
transform -1 0 624 0 1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_41
timestamp -19799
transform -1 0 624 0 -1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_42
timestamp -19799
transform -1 0 624 0 1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_43
timestamp -19799
transform -1 0 624 0 -1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_44
timestamp -19799
transform -1 0 624 0 1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_45
timestamp -19799
transform -1 0 624 0 -1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_46
timestamp -19799
transform -1 0 624 0 1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_47
timestamp -19799
transform -1 0 624 0 -1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_48
timestamp -19799
transform -1 0 624 0 1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_49
timestamp -19799
transform -1 0 624 0 -1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_50
timestamp -19799
transform -1 0 624 0 1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_51
timestamp -19799
transform -1 0 624 0 -1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_52
timestamp -19799
transform -1 0 624 0 1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_53
timestamp -19799
transform -1 0 624 0 -1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_54
timestamp -19799
transform -1 0 624 0 1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_55
timestamp -19799
transform -1 0 624 0 -1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_56
timestamp -19799
transform -1 0 624 0 1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_57
timestamp -19799
transform -1 0 624 0 -1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_58
timestamp -19799
transform -1 0 624 0 1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_59
timestamp -19799
transform -1 0 624 0 -1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_60
timestamp -19799
transform -1 0 624 0 1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_61
timestamp -19799
transform -1 0 624 0 -1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_62
timestamp -19799
transform -1 0 624 0 1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_63
timestamp -19799
transform -1 0 624 0 -1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_64
timestamp -19799
transform -1 0 624 0 1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_65
timestamp -19799
transform -1 0 624 0 -1 790
box -42 -55 624 371
<< labels >>
rlabel metal2 s 0 1113 28 1161 4 wl0_1
port 3 nsew
rlabel metal2 s 0 893 28 941 4 wl1_1
port 5 nsew
rlabel metal2 s 0 1209 28 1257 4 wl0_2
port 7 nsew
rlabel metal2 s 0 1429 28 1477 4 wl1_2
port 9 nsew
rlabel metal2 s 0 1903 28 1951 4 wl0_3
port 11 nsew
rlabel metal2 s 0 1683 28 1731 4 wl1_3
port 13 nsew
rlabel metal2 s 0 1999 28 2047 4 wl0_4
port 15 nsew
rlabel metal2 s 0 2219 28 2267 4 wl1_4
port 17 nsew
rlabel metal2 s 0 2693 28 2741 4 wl0_5
port 19 nsew
rlabel metal2 s 0 2473 28 2521 4 wl1_5
port 21 nsew
rlabel metal2 s 0 2789 28 2837 4 wl0_6
port 23 nsew
rlabel metal2 s 0 3009 28 3057 4 wl1_6
port 25 nsew
rlabel metal2 s 0 3483 28 3531 4 wl0_7
port 27 nsew
rlabel metal2 s 0 3263 28 3311 4 wl1_7
port 29 nsew
rlabel metal2 s 0 3579 28 3627 4 wl0_8
port 31 nsew
rlabel metal2 s 0 3799 28 3847 4 wl1_8
port 33 nsew
rlabel metal2 s 0 4273 28 4321 4 wl0_9
port 35 nsew
rlabel metal2 s 0 4053 28 4101 4 wl1_9
port 37 nsew
rlabel metal2 s 0 4369 28 4417 4 wl0_10
port 39 nsew
rlabel metal2 s 0 4589 28 4637 4 wl1_10
port 41 nsew
rlabel metal2 s 0 5063 28 5111 4 wl0_11
port 43 nsew
rlabel metal2 s 0 4843 28 4891 4 wl1_11
port 45 nsew
rlabel metal2 s 0 5159 28 5207 4 wl0_12
port 47 nsew
rlabel metal2 s 0 5379 28 5427 4 wl1_12
port 49 nsew
rlabel metal2 s 0 5853 28 5901 4 wl0_13
port 51 nsew
rlabel metal2 s 0 5633 28 5681 4 wl1_13
port 53 nsew
rlabel metal2 s 0 5949 28 5997 4 wl0_14
port 55 nsew
rlabel metal2 s 0 6169 28 6217 4 wl1_14
port 57 nsew
rlabel metal2 s 0 6643 28 6691 4 wl0_15
port 59 nsew
rlabel metal2 s 0 6423 28 6471 4 wl1_15
port 61 nsew
rlabel metal2 s 0 6739 28 6787 4 wl0_16
port 63 nsew
rlabel metal2 s 0 6959 28 7007 4 wl1_16
port 65 nsew
rlabel metal2 s 0 7433 28 7481 4 wl0_17
port 67 nsew
rlabel metal2 s 0 7213 28 7261 4 wl1_17
port 69 nsew
rlabel metal2 s 0 7529 28 7577 4 wl0_18
port 71 nsew
rlabel metal2 s 0 7749 28 7797 4 wl1_18
port 73 nsew
rlabel metal2 s 0 8223 28 8271 4 wl0_19
port 75 nsew
rlabel metal2 s 0 8003 28 8051 4 wl1_19
port 77 nsew
rlabel metal2 s 0 8319 28 8367 4 wl0_20
port 79 nsew
rlabel metal2 s 0 8539 28 8587 4 wl1_20
port 81 nsew
rlabel metal2 s 0 9013 28 9061 4 wl0_21
port 83 nsew
rlabel metal2 s 0 8793 28 8841 4 wl1_21
port 85 nsew
rlabel metal2 s 0 9109 28 9157 4 wl0_22
port 87 nsew
rlabel metal2 s 0 9329 28 9377 4 wl1_22
port 89 nsew
rlabel metal2 s 0 9803 28 9851 4 wl0_23
port 91 nsew
rlabel metal2 s 0 9583 28 9631 4 wl1_23
port 93 nsew
rlabel metal2 s 0 9899 28 9947 4 wl0_24
port 95 nsew
rlabel metal2 s 0 10119 28 10167 4 wl1_24
port 97 nsew
rlabel metal2 s 0 10593 28 10641 4 wl0_25
port 99 nsew
rlabel metal2 s 0 10373 28 10421 4 wl1_25
port 101 nsew
rlabel metal2 s 0 10689 28 10737 4 wl0_26
port 103 nsew
rlabel metal2 s 0 10909 28 10957 4 wl1_26
port 105 nsew
rlabel metal2 s 0 11383 28 11431 4 wl0_27
port 107 nsew
rlabel metal2 s 0 11163 28 11211 4 wl1_27
port 109 nsew
rlabel metal2 s 0 11479 28 11527 4 wl0_28
port 111 nsew
rlabel metal2 s 0 11699 28 11747 4 wl1_28
port 113 nsew
rlabel metal2 s 0 12173 28 12221 4 wl0_29
port 115 nsew
rlabel metal2 s 0 11953 28 12001 4 wl1_29
port 117 nsew
rlabel metal2 s 0 12269 28 12317 4 wl0_30
port 119 nsew
rlabel metal2 s 0 12489 28 12537 4 wl1_30
port 121 nsew
rlabel metal2 s 0 12963 28 13011 4 wl0_31
port 123 nsew
rlabel metal2 s 0 12743 28 12791 4 wl1_31
port 125 nsew
rlabel metal2 s 0 13059 28 13107 4 wl0_32
port 127 nsew
rlabel metal2 s 0 13279 28 13327 4 wl1_32
port 129 nsew
rlabel metal2 s 0 13753 28 13801 4 wl0_33
port 131 nsew
rlabel metal2 s 0 13533 28 13581 4 wl1_33
port 133 nsew
rlabel metal2 s 0 13849 28 13897 4 wl0_34
port 135 nsew
rlabel metal2 s 0 14069 28 14117 4 wl1_34
port 137 nsew
rlabel metal2 s 0 14543 28 14591 4 wl0_35
port 139 nsew
rlabel metal2 s 0 14323 28 14371 4 wl1_35
port 141 nsew
rlabel metal2 s 0 14639 28 14687 4 wl0_36
port 143 nsew
rlabel metal2 s 0 14859 28 14907 4 wl1_36
port 145 nsew
rlabel metal2 s 0 15333 28 15381 4 wl0_37
port 147 nsew
rlabel metal2 s 0 15113 28 15161 4 wl1_37
port 149 nsew
rlabel metal2 s 0 15429 28 15477 4 wl0_38
port 151 nsew
rlabel metal2 s 0 15649 28 15697 4 wl1_38
port 153 nsew
rlabel metal2 s 0 16123 28 16171 4 wl0_39
port 155 nsew
rlabel metal2 s 0 15903 28 15951 4 wl1_39
port 157 nsew
rlabel metal2 s 0 16219 28 16267 4 wl0_40
port 159 nsew
rlabel metal2 s 0 16439 28 16487 4 wl1_40
port 161 nsew
rlabel metal2 s 0 16913 28 16961 4 wl0_41
port 163 nsew
rlabel metal2 s 0 16693 28 16741 4 wl1_41
port 165 nsew
rlabel metal2 s 0 17009 28 17057 4 wl0_42
port 167 nsew
rlabel metal2 s 0 17229 28 17277 4 wl1_42
port 169 nsew
rlabel metal2 s 0 17703 28 17751 4 wl0_43
port 171 nsew
rlabel metal2 s 0 17483 28 17531 4 wl1_43
port 173 nsew
rlabel metal2 s 0 17799 28 17847 4 wl0_44
port 175 nsew
rlabel metal2 s 0 18019 28 18067 4 wl1_44
port 177 nsew
rlabel metal2 s 0 18493 28 18541 4 wl0_45
port 179 nsew
rlabel metal2 s 0 18273 28 18321 4 wl1_45
port 181 nsew
rlabel metal2 s 0 18589 28 18637 4 wl0_46
port 183 nsew
rlabel metal2 s 0 18809 28 18857 4 wl1_46
port 185 nsew
rlabel metal2 s 0 19283 28 19331 4 wl0_47
port 187 nsew
rlabel metal2 s 0 19063 28 19111 4 wl1_47
port 189 nsew
rlabel metal2 s 0 19379 28 19427 4 wl0_48
port 191 nsew
rlabel metal2 s 0 19599 28 19647 4 wl1_48
port 193 nsew
rlabel metal2 s 0 20073 28 20121 4 wl0_49
port 195 nsew
rlabel metal2 s 0 19853 28 19901 4 wl1_49
port 197 nsew
rlabel metal2 s 0 20169 28 20217 4 wl0_50
port 199 nsew
rlabel metal2 s 0 20389 28 20437 4 wl1_50
port 201 nsew
rlabel metal2 s 0 20863 28 20911 4 wl0_51
port 203 nsew
rlabel metal2 s 0 20643 28 20691 4 wl1_51
port 205 nsew
rlabel metal2 s 0 20959 28 21007 4 wl0_52
port 207 nsew
rlabel metal2 s 0 21179 28 21227 4 wl1_52
port 209 nsew
rlabel metal2 s 0 21653 28 21701 4 wl0_53
port 211 nsew
rlabel metal2 s 0 21433 28 21481 4 wl1_53
port 213 nsew
rlabel metal2 s 0 21749 28 21797 4 wl0_54
port 215 nsew
rlabel metal2 s 0 21969 28 22017 4 wl1_54
port 217 nsew
rlabel metal2 s 0 22443 28 22491 4 wl0_55
port 219 nsew
rlabel metal2 s 0 22223 28 22271 4 wl1_55
port 221 nsew
rlabel metal2 s 0 22539 28 22587 4 wl0_56
port 223 nsew
rlabel metal2 s 0 22759 28 22807 4 wl1_56
port 225 nsew
rlabel metal2 s 0 23233 28 23281 4 wl0_57
port 227 nsew
rlabel metal2 s 0 23013 28 23061 4 wl1_57
port 229 nsew
rlabel metal2 s 0 23329 28 23377 4 wl0_58
port 231 nsew
rlabel metal2 s 0 23549 28 23597 4 wl1_58
port 233 nsew
rlabel metal2 s 0 24023 28 24071 4 wl0_59
port 235 nsew
rlabel metal2 s 0 23803 28 23851 4 wl1_59
port 237 nsew
rlabel metal2 s 0 24119 28 24167 4 wl0_60
port 239 nsew
rlabel metal2 s 0 24339 28 24387 4 wl1_60
port 241 nsew
rlabel metal2 s 0 24813 28 24861 4 wl0_61
port 243 nsew
rlabel metal2 s 0 24593 28 24641 4 wl1_61
port 245 nsew
rlabel metal2 s 0 24909 28 24957 4 wl0_62
port 247 nsew
rlabel metal2 s 0 25129 28 25177 4 wl1_62
port 249 nsew
rlabel metal2 s 0 25603 28 25651 4 wl0_63
port 251 nsew
rlabel metal2 s 0 25383 28 25431 4 wl1_63
port 253 nsew
rlabel metal2 s 0 25699 28 25747 4 wl0_64
port 255 nsew
rlabel metal2 s 0 25919 28 25967 4 wl1_64
port 257 nsew
rlabel metal2 s 330 989 438 1065 4 gnd
port 259 nsew
rlabel metal2 s 330 1525 438 1635 4 gnd
port 259 nsew
rlabel metal2 s 330 7845 438 7955 4 gnd
port 259 nsew
rlabel metal2 s 330 10215 438 10325 4 gnd
port 259 nsew
rlabel metal2 s 330 9425 438 9535 4 gnd
port 259 nsew
rlabel metal2 s 330 24215 438 24291 4 gnd
port 259 nsew
rlabel metal2 s 330 23899 438 23975 4 gnd
port 259 nsew
rlabel metal2 s 330 19949 438 20025 4 gnd
port 259 nsew
rlabel metal2 s 330 2315 438 2425 4 gnd
port 259 nsew
rlabel metal2 s 330 14165 438 14275 4 gnd
port 259 nsew
rlabel metal2 s 330 6045 438 6121 4 gnd
port 259 nsew
rlabel metal2 s 330 20265 438 20341 4 gnd
port 259 nsew
rlabel metal2 s 330 4685 438 4795 4 gnd
port 259 nsew
rlabel metal2 s 330 1779 438 1855 4 gnd
port 259 nsew
rlabel metal2 s 330 15745 438 15855 4 gnd
port 259 nsew
rlabel metal2 s 330 9679 438 9755 4 gnd
port 259 nsew
rlabel metal2 s 330 10469 438 10545 4 gnd
port 259 nsew
rlabel metal2 s 330 3895 438 4005 4 gnd
port 259 nsew
rlabel metal2 s 330 19159 438 19235 4 gnd
port 259 nsew
rlabel metal2 s 330 18115 438 18225 4 gnd
port 259 nsew
rlabel metal2 s 330 5255 438 5331 4 gnd
port 259 nsew
rlabel metal2 s 330 13629 438 13705 4 gnd
port 259 nsew
rlabel metal2 s 330 3675 438 3751 4 gnd
port 259 nsew
rlabel metal2 s 330 25795 438 25871 4 gnd
port 259 nsew
rlabel metal2 s 330 9205 438 9281 4 gnd
port 259 nsew
rlabel metal2 s 330 14735 438 14811 4 gnd
port 259 nsew
rlabel metal2 s 330 20485 438 20595 4 gnd
port 259 nsew
rlabel metal2 s 330 1305 438 1381 4 gnd
port 259 nsew
rlabel metal2 s 330 6519 438 6595 4 gnd
port 259 nsew
rlabel metal2 s 330 16789 438 16865 4 gnd
port 259 nsew
rlabel metal2 s 330 8635 438 8745 4 gnd
port 259 nsew
rlabel metal2 s 330 10785 438 10861 4 gnd
port 259 nsew
rlabel metal2 s 330 15209 438 15285 4 gnd
port 259 nsew
rlabel metal2 s 330 23425 438 23501 4 gnd
port 259 nsew
rlabel metal2 s 330 4149 438 4225 4 gnd
port 259 nsew
rlabel metal2 s 330 7625 438 7701 4 gnd
port 259 nsew
rlabel metal2 s 330 735 438 845 4 gnd
port 259 nsew
rlabel metal2 s 330 8415 438 8491 4 gnd
port 259 nsew
rlabel metal2 s 330 2885 438 2961 4 gnd
port 259 nsew
rlabel metal2 s 330 11795 438 11905 4 gnd
port 259 nsew
rlabel metal2 s 330 13155 438 13231 4 gnd
port 259 nsew
rlabel metal2 s 330 16535 438 16645 4 gnd
port 259 nsew
rlabel metal2 s 330 11005 438 11115 4 gnd
port 259 nsew
rlabel metal2 s 330 20739 438 20815 4 gnd
port 259 nsew
rlabel metal2 s 330 19475 438 19551 4 gnd
port 259 nsew
rlabel metal2 s 330 22319 438 22395 4 gnd
port 259 nsew
rlabel metal2 s 330 13375 438 13485 4 gnd
port 259 nsew
rlabel metal2 s 330 21845 438 21921 4 gnd
port 259 nsew
rlabel metal2 s 330 16315 438 16391 4 gnd
port 259 nsew
rlabel metal2 s 330 25225 438 25335 4 gnd
port 259 nsew
rlabel metal2 s 330 11575 438 11651 4 gnd
port 259 nsew
rlabel metal2 s 330 24435 438 24545 4 gnd
port 259 nsew
rlabel metal2 s 330 4465 438 4541 4 gnd
port 259 nsew
rlabel metal2 s 330 25479 438 25555 4 gnd
port 259 nsew
rlabel metal2 s 330 13945 438 14021 4 gnd
port 259 nsew
rlabel metal2 s 330 24689 438 24765 4 gnd
port 259 nsew
rlabel metal2 s 330 14955 438 15065 4 gnd
port 259 nsew
rlabel metal2 s 330 17325 438 17435 4 gnd
port 259 nsew
rlabel metal2 s 330 6835 438 6911 4 gnd
port 259 nsew
rlabel metal2 s 330 3105 438 3215 4 gnd
port 259 nsew
rlabel metal2 s 330 5475 438 5585 4 gnd
port 259 nsew
rlabel metal2 s 330 23645 438 23755 4 gnd
port 259 nsew
rlabel metal2 s 330 9995 438 10071 4 gnd
port 259 nsew
rlabel metal2 s 330 18369 438 18445 4 gnd
port 259 nsew
rlabel metal2 s 330 8099 438 8175 4 gnd
port 259 nsew
rlabel metal2 s 330 2095 438 2171 4 gnd
port 259 nsew
rlabel metal2 s 330 3359 438 3435 4 gnd
port 259 nsew
rlabel metal2 s 330 22635 438 22711 4 gnd
port 259 nsew
rlabel metal2 s 330 22065 438 22175 4 gnd
port 259 nsew
rlabel metal2 s 330 17895 438 17971 4 gnd
port 259 nsew
rlabel metal2 s 330 23109 438 23185 4 gnd
port 259 nsew
rlabel metal2 s 330 11259 438 11335 4 gnd
port 259 nsew
rlabel metal2 s 330 15525 438 15601 4 gnd
port 259 nsew
rlabel metal2 s 330 18905 438 19015 4 gnd
port 259 nsew
rlabel metal2 s 330 25005 438 25081 4 gnd
port 259 nsew
rlabel metal2 s 330 12365 438 12441 4 gnd
port 259 nsew
rlabel metal2 s 330 4939 438 5015 4 gnd
port 259 nsew
rlabel metal2 s 330 18685 438 18761 4 gnd
port 259 nsew
rlabel metal2 s 330 17105 438 17181 4 gnd
port 259 nsew
rlabel metal2 s 330 6265 438 6375 4 gnd
port 259 nsew
rlabel metal2 s 330 15999 438 16075 4 gnd
port 259 nsew
rlabel metal2 s 330 21055 438 21131 4 gnd
port 259 nsew
rlabel metal2 s 330 14419 438 14495 4 gnd
port 259 nsew
rlabel metal2 s 330 21529 438 21605 4 gnd
port 259 nsew
rlabel metal2 s 330 21275 438 21385 4 gnd
port 259 nsew
rlabel metal2 s 330 2569 438 2645 4 gnd
port 259 nsew
rlabel metal2 s 330 22855 438 22965 4 gnd
port 259 nsew
rlabel metal2 s 330 7055 438 7165 4 gnd
port 259 nsew
rlabel metal2 s 330 12049 438 12125 4 gnd
port 259 nsew
rlabel metal2 s 330 8889 438 8965 4 gnd
port 259 nsew
rlabel metal2 s 330 7309 438 7385 4 gnd
port 259 nsew
rlabel metal2 s 330 5729 438 5805 4 gnd
port 259 nsew
rlabel metal2 s 330 12585 438 12695 4 gnd
port 259 nsew
rlabel metal2 s 330 26015 438 26125 4 gnd
port 259 nsew
rlabel metal2 s 330 12839 438 12915 4 gnd
port 259 nsew
rlabel metal2 s 330 19695 438 19805 4 gnd
port 259 nsew
rlabel metal2 s 330 17579 438 17655 4 gnd
port 259 nsew
<< properties >>
string FIXED_BBOX 0 0 624 26465
<< end >>
