magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1195 -1260 1935 2576
<< pwell >>
rect 211 730 413 1286
rect 211 596 675 730
rect 211 28 413 596
<< scnmos >>
rect 297 684 327 1260
rect 297 54 327 630
<< ndiff >>
rect 237 989 297 1260
rect 237 955 245 989
rect 279 955 297 989
rect 237 684 297 955
rect 327 989 387 1260
rect 327 955 345 989
rect 379 955 387 989
rect 327 684 387 955
rect 237 359 297 630
rect 237 325 245 359
rect 279 325 297 359
rect 237 54 297 325
rect 327 359 387 630
rect 327 325 345 359
rect 379 325 387 359
rect 327 54 387 325
<< ndiffc >>
rect 245 955 279 989
rect 345 955 379 989
rect 245 325 279 359
rect 345 325 379 359
<< psubdiff >>
rect 599 680 649 704
rect 599 646 607 680
rect 641 646 649 680
rect 599 622 649 646
<< psubdiffcont >>
rect 607 646 641 680
<< poly >>
rect 297 1260 327 1286
rect 297 630 327 684
rect 297 28 327 54
<< locali >>
rect 77 1277 111 1293
rect 111 1243 379 1277
rect 77 1227 111 1243
rect 245 989 279 1005
rect 245 939 279 955
rect 345 989 379 1243
rect 345 939 379 955
rect 607 680 641 696
rect 607 630 641 646
rect 245 359 279 375
rect 245 73 279 325
rect 345 359 379 375
rect 345 309 379 325
rect 541 73 575 89
rect 245 39 541 73
rect 541 23 575 39
<< viali >>
rect 77 1243 111 1277
rect 245 955 279 989
rect 607 646 641 680
rect 345 325 379 359
rect 541 39 575 73
<< metal1 >>
rect 80 1283 108 1316
rect 65 1277 123 1283
rect 65 1243 77 1277
rect 111 1243 123 1277
rect 65 1237 123 1243
rect 233 989 291 995
rect 233 955 245 989
rect 279 955 291 989
rect 233 949 291 955
rect 248 412 276 949
rect 544 832 572 1316
rect 80 384 276 412
rect 348 804 572 832
rect 80 0 108 384
rect 348 365 376 804
rect 595 680 653 686
rect 595 646 607 680
rect 641 646 653 680
rect 595 640 653 646
rect 333 359 391 365
rect 333 325 345 359
rect 379 325 391 359
rect 333 319 391 325
rect 529 73 587 79
rect 529 39 541 73
rect 575 39 587 73
rect 529 33 587 39
rect 544 0 572 33
<< labels >>
rlabel poly s 312 41 312 41 4 sel
port 2 nsew
rlabel metal1 s 80 1260 108 1316 4 bl
port 4 nsew
rlabel metal1 s 544 1260 572 1316 4 br
port 6 nsew
rlabel metal1 s 80 0 108 56 4 bl_out
port 8 nsew
rlabel metal1 s 544 0 572 56 4 br_out
port 10 nsew
rlabel metal1 s 610 649 638 677 4 gnd
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 624 597
<< end >>
