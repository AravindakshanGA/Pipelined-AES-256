magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1260 -1008 23180 6929
<< metal1 >>
rect 2142 5613 2202 5669
rect 4638 5613 4698 5669
rect 7134 5613 7194 5669
rect 9630 5613 9690 5669
rect 12126 5613 12186 5669
rect 14622 5613 14682 5669
rect 17118 5613 17178 5669
rect 19614 5613 19674 5669
rect 0 5551 19891 5579
rect 2046 3596 2074 3662
rect 1999 3568 2074 3596
rect 1999 3162 2027 3568
rect 2248 3516 2276 3662
rect 4542 3596 4570 3662
rect 4495 3568 4570 3596
rect 2248 3488 2491 3516
rect 2463 3286 2491 3488
rect 4495 3162 4523 3568
rect 4744 3516 4772 3662
rect 7038 3596 7066 3662
rect 6991 3568 7066 3596
rect 4744 3488 4987 3516
rect 4959 3286 4987 3488
rect 6991 3162 7019 3568
rect 7240 3516 7268 3662
rect 9534 3596 9562 3662
rect 9487 3568 9562 3596
rect 7240 3488 7483 3516
rect 7455 3286 7483 3488
rect 9487 3162 9515 3568
rect 9736 3516 9764 3662
rect 12030 3596 12058 3662
rect 11983 3568 12058 3596
rect 9736 3488 9979 3516
rect 9951 3286 9979 3488
rect 11983 3162 12011 3568
rect 12232 3516 12260 3662
rect 14526 3596 14554 3662
rect 14479 3568 14554 3596
rect 12232 3488 12475 3516
rect 12447 3286 12475 3488
rect 14479 3162 14507 3568
rect 14728 3516 14756 3662
rect 17022 3596 17050 3662
rect 16975 3568 17050 3596
rect 14728 3488 14971 3516
rect 14943 3286 14971 3488
rect 16975 3162 17003 3568
rect 17224 3516 17252 3662
rect 19518 3596 19546 3662
rect 19471 3568 19546 3596
rect 17224 3488 17467 3516
rect 17439 3286 17467 3488
rect 19471 3162 19499 3568
rect 19720 3516 19748 3662
rect 19720 3488 19963 3516
rect 19935 3286 19963 3488
rect 1999 1160 2027 1226
rect 1985 1132 2027 1160
rect 1361 252 1389 974
rect 1825 252 1853 974
rect 1985 252 2013 1132
rect 2463 1080 2491 1226
rect 2449 1052 2491 1080
rect 2595 1080 2623 1226
rect 3059 1160 3087 1226
rect 3247 1160 3275 1226
rect 3059 1132 3101 1160
rect 2595 1052 2637 1080
rect 2449 252 2477 1052
rect 2609 252 2637 1052
rect 3073 252 3101 1132
rect 3233 1132 3275 1160
rect 3233 252 3261 1132
rect 3711 1080 3739 1226
rect 3697 1052 3739 1080
rect 3843 1080 3871 1226
rect 4307 1160 4335 1226
rect 4495 1160 4523 1226
rect 4307 1132 4349 1160
rect 3843 1052 3885 1080
rect 3697 252 3725 1052
rect 3857 252 3885 1052
rect 4321 252 4349 1132
rect 4481 1132 4523 1160
rect 4481 252 4509 1132
rect 4959 1080 4987 1226
rect 4945 1052 4987 1080
rect 5091 1080 5119 1226
rect 5555 1160 5583 1226
rect 5743 1160 5771 1226
rect 5555 1132 5597 1160
rect 5091 1052 5133 1080
rect 4945 252 4973 1052
rect 5105 252 5133 1052
rect 5569 252 5597 1132
rect 5729 1132 5771 1160
rect 5729 252 5757 1132
rect 6207 1080 6235 1226
rect 6193 1052 6235 1080
rect 6339 1080 6367 1226
rect 6803 1160 6831 1226
rect 6991 1160 7019 1226
rect 6803 1132 6845 1160
rect 6339 1052 6381 1080
rect 6193 252 6221 1052
rect 6353 252 6381 1052
rect 6817 252 6845 1132
rect 6977 1132 7019 1160
rect 6977 252 7005 1132
rect 7455 1080 7483 1226
rect 7441 1052 7483 1080
rect 7587 1080 7615 1226
rect 8051 1160 8079 1226
rect 8239 1160 8267 1226
rect 8051 1132 8093 1160
rect 7587 1052 7629 1080
rect 7441 252 7469 1052
rect 7601 252 7629 1052
rect 8065 252 8093 1132
rect 8225 1132 8267 1160
rect 8225 252 8253 1132
rect 8703 1080 8731 1226
rect 8689 1052 8731 1080
rect 8835 1080 8863 1226
rect 9299 1160 9327 1226
rect 9487 1160 9515 1226
rect 9299 1132 9341 1160
rect 8835 1052 8877 1080
rect 8689 252 8717 1052
rect 8849 252 8877 1052
rect 9313 252 9341 1132
rect 9473 1132 9515 1160
rect 9473 252 9501 1132
rect 9951 1080 9979 1226
rect 9937 1052 9979 1080
rect 10083 1080 10111 1226
rect 10547 1160 10575 1226
rect 10735 1160 10763 1226
rect 10547 1132 10589 1160
rect 10083 1052 10125 1080
rect 9937 252 9965 1052
rect 10097 252 10125 1052
rect 10561 252 10589 1132
rect 10721 1132 10763 1160
rect 10721 252 10749 1132
rect 11199 1080 11227 1226
rect 11185 1052 11227 1080
rect 11331 1080 11359 1226
rect 11795 1160 11823 1226
rect 11983 1160 12011 1226
rect 11795 1132 11837 1160
rect 11331 1052 11373 1080
rect 11185 252 11213 1052
rect 11345 252 11373 1052
rect 11809 252 11837 1132
rect 11969 1132 12011 1160
rect 11969 252 11997 1132
rect 12447 1080 12475 1226
rect 12433 1052 12475 1080
rect 12579 1080 12607 1226
rect 13043 1160 13071 1226
rect 13231 1160 13259 1226
rect 13043 1132 13085 1160
rect 12579 1052 12621 1080
rect 12433 252 12461 1052
rect 12593 252 12621 1052
rect 13057 252 13085 1132
rect 13217 1132 13259 1160
rect 13217 252 13245 1132
rect 13695 1080 13723 1226
rect 13681 1052 13723 1080
rect 13827 1080 13855 1226
rect 14291 1160 14319 1226
rect 14479 1160 14507 1226
rect 14291 1132 14333 1160
rect 13827 1052 13869 1080
rect 13681 252 13709 1052
rect 13841 252 13869 1052
rect 14305 252 14333 1132
rect 14465 1132 14507 1160
rect 14465 252 14493 1132
rect 14943 1080 14971 1226
rect 14929 1052 14971 1080
rect 15075 1080 15103 1226
rect 15539 1160 15567 1226
rect 15727 1160 15755 1226
rect 15539 1132 15581 1160
rect 15075 1052 15117 1080
rect 14929 252 14957 1052
rect 15089 252 15117 1052
rect 15553 252 15581 1132
rect 15713 1132 15755 1160
rect 15713 252 15741 1132
rect 16191 1080 16219 1226
rect 16177 1052 16219 1080
rect 16323 1080 16351 1226
rect 16787 1160 16815 1226
rect 16975 1160 17003 1226
rect 16787 1132 16829 1160
rect 16323 1052 16365 1080
rect 16177 252 16205 1052
rect 16337 252 16365 1052
rect 16801 252 16829 1132
rect 16961 1132 17003 1160
rect 16961 252 16989 1132
rect 17439 1080 17467 1226
rect 17425 1052 17467 1080
rect 17571 1080 17599 1226
rect 18035 1160 18063 1226
rect 18223 1160 18251 1226
rect 18035 1132 18077 1160
rect 17571 1052 17613 1080
rect 17425 252 17453 1052
rect 17585 252 17613 1052
rect 18049 252 18077 1132
rect 18209 1132 18251 1160
rect 18209 252 18237 1132
rect 18687 1080 18715 1226
rect 18673 1052 18715 1080
rect 18819 1080 18847 1226
rect 19283 1160 19311 1226
rect 19471 1160 19499 1226
rect 19283 1132 19325 1160
rect 18819 1052 18861 1080
rect 18673 252 18701 1052
rect 18833 252 18861 1052
rect 19297 252 19325 1132
rect 19457 1132 19499 1160
rect 19457 252 19485 1132
rect 19935 1080 19963 1226
rect 19921 1052 19963 1080
rect 20067 1080 20095 1226
rect 20531 1160 20559 1226
rect 20719 1160 20747 1226
rect 20531 1132 20573 1160
rect 20067 1052 20109 1080
rect 19921 252 19949 1052
rect 20081 252 20109 1052
rect 20545 252 20573 1132
rect 20705 1132 20747 1160
rect 20705 252 20733 1132
rect 21183 1080 21211 1226
rect 21169 1052 21211 1080
rect 21315 1080 21343 1226
rect 21779 1160 21807 1226
rect 21779 1132 21821 1160
rect 21315 1052 21357 1080
rect 21169 252 21197 1052
rect 21329 252 21357 1052
rect 21793 252 21821 1132
<< metal3 >>
rect 33 5323 19924 5389
rect 33 4831 19924 4897
rect 33 4499 19924 4565
rect 33 4062 19924 4128
rect 0 2978 21887 3038
rect 0 2854 21887 2914
rect 0 2730 21887 2790
rect 0 2606 21887 2666
rect 33 1846 21310 1912
rect 33 916 21920 982
rect 33 313 21920 379
use subbyte2_column_mux_array  subbyte2_column_mux_array_0
timestamp 1543373570
transform 1 0 0 0 -1 3410
box 0 87 21887 2184
use subbyte2_precharge_array  subbyte2_precharge_array_0
timestamp 1543373570
transform 1 0 0 0 -1 974
box 33 -12 21920 722
use subbyte2_write_driver_array  subbyte2_write_driver_array_0
timestamp 1543373570
transform 1 0 0 0 -1 5673
box 0 4 20271 2011
<< labels >>
rlabel metal1 s 2142 5613 2202 5669 4 din_0
port 3 nsew
rlabel metal1 s 4638 5613 4698 5669 4 din_1
port 5 nsew
rlabel metal1 s 7134 5613 7194 5669 4 din_2
port 7 nsew
rlabel metal1 s 9630 5613 9690 5669 4 din_3
port 9 nsew
rlabel metal1 s 12126 5613 12186 5669 4 din_4
port 11 nsew
rlabel metal1 s 14622 5613 14682 5669 4 din_5
port 13 nsew
rlabel metal1 s 17118 5613 17178 5669 4 din_6
port 15 nsew
rlabel metal1 s 19614 5613 19674 5669 4 din_7
port 17 nsew
rlabel metal1 s 1825 252 1853 974 4 rbl_bl
port 19 nsew
rlabel metal1 s 1361 252 1389 974 4 rbl_br
port 21 nsew
rlabel metal1 s 1985 252 2013 974 4 bl_0
port 23 nsew
rlabel metal1 s 2449 252 2477 974 4 br_0
port 25 nsew
rlabel metal1 s 3073 252 3101 974 4 bl_1
port 27 nsew
rlabel metal1 s 2609 252 2637 974 4 br_1
port 29 nsew
rlabel metal1 s 3233 252 3261 974 4 bl_2
port 31 nsew
rlabel metal1 s 3697 252 3725 974 4 br_2
port 33 nsew
rlabel metal1 s 4321 252 4349 974 4 bl_3
port 35 nsew
rlabel metal1 s 3857 252 3885 974 4 br_3
port 37 nsew
rlabel metal1 s 4481 252 4509 974 4 bl_4
port 39 nsew
rlabel metal1 s 4945 252 4973 974 4 br_4
port 41 nsew
rlabel metal1 s 5569 252 5597 974 4 bl_5
port 43 nsew
rlabel metal1 s 5105 252 5133 974 4 br_5
port 45 nsew
rlabel metal1 s 5729 252 5757 974 4 bl_6
port 47 nsew
rlabel metal1 s 6193 252 6221 974 4 br_6
port 49 nsew
rlabel metal1 s 6817 252 6845 974 4 bl_7
port 51 nsew
rlabel metal1 s 6353 252 6381 974 4 br_7
port 53 nsew
rlabel metal1 s 6977 252 7005 974 4 bl_8
port 55 nsew
rlabel metal1 s 7441 252 7469 974 4 br_8
port 57 nsew
rlabel metal1 s 8065 252 8093 974 4 bl_9
port 59 nsew
rlabel metal1 s 7601 252 7629 974 4 br_9
port 61 nsew
rlabel metal1 s 8225 252 8253 974 4 bl_10
port 63 nsew
rlabel metal1 s 8689 252 8717 974 4 br_10
port 65 nsew
rlabel metal1 s 9313 252 9341 974 4 bl_11
port 67 nsew
rlabel metal1 s 8849 252 8877 974 4 br_11
port 69 nsew
rlabel metal1 s 9473 252 9501 974 4 bl_12
port 71 nsew
rlabel metal1 s 9937 252 9965 974 4 br_12
port 73 nsew
rlabel metal1 s 10561 252 10589 974 4 bl_13
port 75 nsew
rlabel metal1 s 10097 252 10125 974 4 br_13
port 77 nsew
rlabel metal1 s 10721 252 10749 974 4 bl_14
port 79 nsew
rlabel metal1 s 11185 252 11213 974 4 br_14
port 81 nsew
rlabel metal1 s 11809 252 11837 974 4 bl_15
port 83 nsew
rlabel metal1 s 11345 252 11373 974 4 br_15
port 85 nsew
rlabel metal1 s 11969 252 11997 974 4 bl_16
port 87 nsew
rlabel metal1 s 12433 252 12461 974 4 br_16
port 89 nsew
rlabel metal1 s 13057 252 13085 974 4 bl_17
port 91 nsew
rlabel metal1 s 12593 252 12621 974 4 br_17
port 93 nsew
rlabel metal1 s 13217 252 13245 974 4 bl_18
port 95 nsew
rlabel metal1 s 13681 252 13709 974 4 br_18
port 97 nsew
rlabel metal1 s 14305 252 14333 974 4 bl_19
port 99 nsew
rlabel metal1 s 13841 252 13869 974 4 br_19
port 101 nsew
rlabel metal1 s 14465 252 14493 974 4 bl_20
port 103 nsew
rlabel metal1 s 14929 252 14957 974 4 br_20
port 105 nsew
rlabel metal1 s 15553 252 15581 974 4 bl_21
port 107 nsew
rlabel metal1 s 15089 252 15117 974 4 br_21
port 109 nsew
rlabel metal1 s 15713 252 15741 974 4 bl_22
port 111 nsew
rlabel metal1 s 16177 252 16205 974 4 br_22
port 113 nsew
rlabel metal1 s 16801 252 16829 974 4 bl_23
port 115 nsew
rlabel metal1 s 16337 252 16365 974 4 br_23
port 117 nsew
rlabel metal1 s 16961 252 16989 974 4 bl_24
port 119 nsew
rlabel metal1 s 17425 252 17453 974 4 br_24
port 121 nsew
rlabel metal1 s 18049 252 18077 974 4 bl_25
port 123 nsew
rlabel metal1 s 17585 252 17613 974 4 br_25
port 125 nsew
rlabel metal1 s 18209 252 18237 974 4 bl_26
port 127 nsew
rlabel metal1 s 18673 252 18701 974 4 br_26
port 129 nsew
rlabel metal1 s 19297 252 19325 974 4 bl_27
port 131 nsew
rlabel metal1 s 18833 252 18861 974 4 br_27
port 133 nsew
rlabel metal1 s 19457 252 19485 974 4 bl_28
port 135 nsew
rlabel metal1 s 19921 252 19949 974 4 br_28
port 137 nsew
rlabel metal1 s 20545 252 20573 974 4 bl_29
port 139 nsew
rlabel metal1 s 20081 252 20109 974 4 br_29
port 141 nsew
rlabel metal1 s 20705 252 20733 974 4 bl_30
port 143 nsew
rlabel metal1 s 21169 252 21197 974 4 br_30
port 145 nsew
rlabel metal1 s 21793 252 21821 974 4 bl_31
port 147 nsew
rlabel metal1 s 21329 252 21357 974 4 br_31
port 149 nsew
rlabel metal3 s 33 916 21920 982 4 p_en_bar
port 151 nsew
rlabel metal3 s 0 2978 21887 3038 4 sel_0
port 153 nsew
rlabel metal3 s 0 2854 21887 2914 4 sel_1
port 155 nsew
rlabel metal3 s 0 2730 21887 2790 4 sel_2
port 157 nsew
rlabel metal3 s 0 2606 21887 2666 4 sel_3
port 159 nsew
rlabel metal1 s 0 5551 19891 5579 4 w_en
port 161 nsew
rlabel metal3 s 33 313 21920 379 4 vdd
port 163 nsew
rlabel metal3 s 33 5323 19924 5389 4 vdd
port 163 nsew
rlabel metal3 s 33 4499 19924 4565 4 vdd
port 163 nsew
rlabel metal3 s 33 4831 19924 4897 4 gnd
port 165 nsew
rlabel metal3 s 33 4062 19924 4128 4 gnd
port 165 nsew
rlabel metal3 s 33 1846 21310 1912 4 gnd
port 165 nsew
<< properties >>
string FIXED_BBOX 0 0 21887 5673
<< end >>
