magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1260 -1260 21588 3816
<< metal1 >>
rect 2010 2468 2016 2520
rect 2068 2468 2074 2520
rect 2115 1430 2149 2556
rect 2191 1442 2219 2556
rect 4506 2468 4512 2520
rect 4564 2468 4570 2520
rect 2338 2316 2344 2368
rect 2396 2316 2402 2368
rect 2256 1542 2262 1594
rect 2314 1542 2320 1594
rect 4611 1430 4645 2556
rect 4687 1442 4715 2556
rect 7002 2468 7008 2520
rect 7060 2468 7066 2520
rect 4834 2316 4840 2368
rect 4892 2316 4898 2368
rect 4752 1542 4758 1594
rect 4810 1542 4816 1594
rect 7107 1430 7141 2556
rect 7183 1442 7211 2556
rect 9498 2468 9504 2520
rect 9556 2468 9562 2520
rect 7330 2316 7336 2368
rect 7388 2316 7394 2368
rect 7248 1542 7254 1594
rect 7306 1542 7312 1594
rect 9603 1430 9637 2556
rect 9679 1442 9707 2556
rect 11994 2468 12000 2520
rect 12052 2468 12058 2520
rect 9826 2316 9832 2368
rect 9884 2316 9890 2368
rect 9744 1542 9750 1594
rect 9802 1542 9808 1594
rect 12099 1430 12133 2556
rect 12175 1442 12203 2556
rect 14490 2468 14496 2520
rect 14548 2468 14554 2520
rect 12322 2316 12328 2368
rect 12380 2316 12386 2368
rect 12240 1542 12246 1594
rect 12298 1542 12304 1594
rect 14595 1430 14629 2556
rect 14671 1442 14699 2556
rect 16986 2468 16992 2520
rect 17044 2468 17050 2520
rect 14818 2316 14824 2368
rect 14876 2316 14882 2368
rect 14736 1542 14742 1594
rect 14794 1542 14800 1594
rect 17091 1430 17125 2556
rect 17167 1442 17195 2556
rect 19482 2468 19488 2520
rect 19540 2468 19546 2520
rect 17314 2316 17320 2368
rect 17372 2316 17378 2368
rect 17232 1542 17238 1594
rect 17290 1542 17296 1594
rect 19587 1430 19621 2556
rect 19663 1442 19691 2556
rect 19810 2316 19816 2368
rect 19868 2316 19874 2368
rect 19728 1542 19734 1594
rect 19786 1542 19792 1594
rect 2268 704 2274 756
rect 2326 704 2332 756
rect 4764 704 4770 756
rect 4822 704 4828 756
rect 7260 704 7266 756
rect 7318 704 7324 756
rect 9756 704 9762 756
rect 9814 704 9820 756
rect 12252 704 12258 756
rect 12310 704 12316 756
rect 14748 704 14754 756
rect 14806 704 14812 756
rect 17244 704 17250 756
rect 17302 704 17308 756
rect 19740 704 19746 756
rect 19798 704 19804 756
rect 2268 382 2274 434
rect 2326 382 2332 434
rect 4764 382 4770 434
rect 4822 382 4828 434
rect 7260 382 7266 434
rect 7318 382 7324 434
rect 9756 382 9762 434
rect 9814 382 9820 434
rect 12252 382 12258 434
rect 12310 382 12316 434
rect 14748 382 14754 434
rect 14806 382 14812 434
rect 17244 382 17250 434
rect 17302 382 17308 434
rect 19740 382 19746 434
rect 19798 382 19804 434
rect 2023 0 2069 150
rect 4519 0 4565 150
rect 7015 0 7061 150
rect 9511 0 9557 150
rect 12007 0 12053 150
rect 14503 0 14549 150
rect 16999 0 17045 150
rect 19495 0 19541 150
<< via1 >>
rect 2016 2468 2068 2520
rect 4512 2468 4564 2520
rect 2344 2316 2396 2368
rect 2262 1542 2314 1594
rect 7008 2468 7060 2520
rect 4840 2316 4892 2368
rect 4758 1542 4810 1594
rect 9504 2468 9556 2520
rect 7336 2316 7388 2368
rect 7254 1542 7306 1594
rect 12000 2468 12052 2520
rect 9832 2316 9884 2368
rect 9750 1542 9802 1594
rect 14496 2468 14548 2520
rect 12328 2316 12380 2368
rect 12246 1542 12298 1594
rect 16992 2468 17044 2520
rect 14824 2316 14876 2368
rect 14742 1542 14794 1594
rect 19488 2468 19540 2520
rect 17320 2316 17372 2368
rect 17238 1542 17290 1594
rect 19816 2316 19868 2368
rect 19734 1542 19786 1594
rect 2274 704 2326 756
rect 4770 704 4822 756
rect 7266 704 7318 756
rect 9762 704 9814 756
rect 12258 704 12310 756
rect 14754 704 14806 756
rect 17250 704 17302 756
rect 19746 704 19798 756
rect 2274 382 2326 434
rect 4770 382 4822 434
rect 7266 382 7318 434
rect 9762 382 9814 434
rect 12258 382 12310 434
rect 14754 382 14806 434
rect 17250 382 17302 434
rect 19746 382 19798 434
<< metal2 >>
rect 2014 2522 2070 2531
rect 2014 2457 2070 2466
rect 4510 2522 4566 2531
rect 4510 2457 4566 2466
rect 7006 2522 7062 2531
rect 7006 2457 7062 2466
rect 9502 2522 9558 2531
rect 9502 2457 9558 2466
rect 11998 2522 12054 2531
rect 11998 2457 12054 2466
rect 14494 2522 14550 2531
rect 14494 2457 14550 2466
rect 16990 2522 17046 2531
rect 16990 2457 17046 2466
rect 19486 2522 19542 2531
rect 19486 2457 19542 2466
rect 2342 2370 2398 2379
rect 2342 2305 2398 2314
rect 4838 2370 4894 2379
rect 4838 2305 4894 2314
rect 7334 2370 7390 2379
rect 7334 2305 7390 2314
rect 9830 2370 9886 2379
rect 9830 2305 9886 2314
rect 12326 2370 12382 2379
rect 12326 2305 12382 2314
rect 14822 2370 14878 2379
rect 14822 2305 14878 2314
rect 17318 2370 17374 2379
rect 17318 2305 17374 2314
rect 19814 2370 19870 2379
rect 19814 2305 19870 2314
rect 2260 1596 2316 1605
rect 2260 1531 2316 1540
rect 4756 1596 4812 1605
rect 4756 1531 4812 1540
rect 7252 1596 7308 1605
rect 7252 1531 7308 1540
rect 9748 1596 9804 1605
rect 9748 1531 9804 1540
rect 12244 1596 12300 1605
rect 12244 1531 12300 1540
rect 14740 1596 14796 1605
rect 14740 1531 14796 1540
rect 17236 1596 17292 1605
rect 17236 1531 17292 1540
rect 19732 1596 19788 1605
rect 19732 1531 19788 1540
rect 2272 758 2328 767
rect 2272 693 2328 702
rect 4768 758 4824 767
rect 4768 693 4824 702
rect 7264 758 7320 767
rect 7264 693 7320 702
rect 9760 758 9816 767
rect 9760 693 9816 702
rect 12256 758 12312 767
rect 12256 693 12312 702
rect 14752 758 14808 767
rect 14752 693 14808 702
rect 17248 758 17304 767
rect 17248 693 17304 702
rect 19744 758 19800 767
rect 19744 693 19800 702
rect 2272 436 2328 445
rect 2272 371 2328 380
rect 4768 436 4824 445
rect 4768 371 4824 380
rect 7264 436 7320 445
rect 7264 371 7320 380
rect 9760 436 9816 445
rect 9760 371 9816 380
rect 12256 436 12312 445
rect 12256 371 12312 380
rect 14752 436 14808 445
rect 14752 371 14808 380
rect 17248 436 17304 445
rect 17248 371 17304 380
rect 19744 436 19800 445
rect 19744 371 19800 380
<< via2 >>
rect 2014 2520 2070 2522
rect 2014 2468 2016 2520
rect 2016 2468 2068 2520
rect 2068 2468 2070 2520
rect 2014 2466 2070 2468
rect 4510 2520 4566 2522
rect 4510 2468 4512 2520
rect 4512 2468 4564 2520
rect 4564 2468 4566 2520
rect 4510 2466 4566 2468
rect 7006 2520 7062 2522
rect 7006 2468 7008 2520
rect 7008 2468 7060 2520
rect 7060 2468 7062 2520
rect 7006 2466 7062 2468
rect 9502 2520 9558 2522
rect 9502 2468 9504 2520
rect 9504 2468 9556 2520
rect 9556 2468 9558 2520
rect 9502 2466 9558 2468
rect 11998 2520 12054 2522
rect 11998 2468 12000 2520
rect 12000 2468 12052 2520
rect 12052 2468 12054 2520
rect 11998 2466 12054 2468
rect 14494 2520 14550 2522
rect 14494 2468 14496 2520
rect 14496 2468 14548 2520
rect 14548 2468 14550 2520
rect 14494 2466 14550 2468
rect 16990 2520 17046 2522
rect 16990 2468 16992 2520
rect 16992 2468 17044 2520
rect 17044 2468 17046 2520
rect 16990 2466 17046 2468
rect 19486 2520 19542 2522
rect 19486 2468 19488 2520
rect 19488 2468 19540 2520
rect 19540 2468 19542 2520
rect 19486 2466 19542 2468
rect 2342 2368 2398 2370
rect 2342 2316 2344 2368
rect 2344 2316 2396 2368
rect 2396 2316 2398 2368
rect 2342 2314 2398 2316
rect 4838 2368 4894 2370
rect 4838 2316 4840 2368
rect 4840 2316 4892 2368
rect 4892 2316 4894 2368
rect 4838 2314 4894 2316
rect 7334 2368 7390 2370
rect 7334 2316 7336 2368
rect 7336 2316 7388 2368
rect 7388 2316 7390 2368
rect 7334 2314 7390 2316
rect 9830 2368 9886 2370
rect 9830 2316 9832 2368
rect 9832 2316 9884 2368
rect 9884 2316 9886 2368
rect 9830 2314 9886 2316
rect 12326 2368 12382 2370
rect 12326 2316 12328 2368
rect 12328 2316 12380 2368
rect 12380 2316 12382 2368
rect 12326 2314 12382 2316
rect 14822 2368 14878 2370
rect 14822 2316 14824 2368
rect 14824 2316 14876 2368
rect 14876 2316 14878 2368
rect 14822 2314 14878 2316
rect 17318 2368 17374 2370
rect 17318 2316 17320 2368
rect 17320 2316 17372 2368
rect 17372 2316 17374 2368
rect 17318 2314 17374 2316
rect 19814 2368 19870 2370
rect 19814 2316 19816 2368
rect 19816 2316 19868 2368
rect 19868 2316 19870 2368
rect 19814 2314 19870 2316
rect 2260 1594 2316 1596
rect 2260 1542 2262 1594
rect 2262 1542 2314 1594
rect 2314 1542 2316 1594
rect 2260 1540 2316 1542
rect 4756 1594 4812 1596
rect 4756 1542 4758 1594
rect 4758 1542 4810 1594
rect 4810 1542 4812 1594
rect 4756 1540 4812 1542
rect 7252 1594 7308 1596
rect 7252 1542 7254 1594
rect 7254 1542 7306 1594
rect 7306 1542 7308 1594
rect 7252 1540 7308 1542
rect 9748 1594 9804 1596
rect 9748 1542 9750 1594
rect 9750 1542 9802 1594
rect 9802 1542 9804 1594
rect 9748 1540 9804 1542
rect 12244 1594 12300 1596
rect 12244 1542 12246 1594
rect 12246 1542 12298 1594
rect 12298 1542 12300 1594
rect 12244 1540 12300 1542
rect 14740 1594 14796 1596
rect 14740 1542 14742 1594
rect 14742 1542 14794 1594
rect 14794 1542 14796 1594
rect 14740 1540 14796 1542
rect 17236 1594 17292 1596
rect 17236 1542 17238 1594
rect 17238 1542 17290 1594
rect 17290 1542 17292 1594
rect 17236 1540 17292 1542
rect 19732 1594 19788 1596
rect 19732 1542 19734 1594
rect 19734 1542 19786 1594
rect 19786 1542 19788 1594
rect 19732 1540 19788 1542
rect 2272 756 2328 758
rect 2272 704 2274 756
rect 2274 704 2326 756
rect 2326 704 2328 756
rect 2272 702 2328 704
rect 4768 756 4824 758
rect 4768 704 4770 756
rect 4770 704 4822 756
rect 4822 704 4824 756
rect 4768 702 4824 704
rect 7264 756 7320 758
rect 7264 704 7266 756
rect 7266 704 7318 756
rect 7318 704 7320 756
rect 7264 702 7320 704
rect 9760 756 9816 758
rect 9760 704 9762 756
rect 9762 704 9814 756
rect 9814 704 9816 756
rect 9760 702 9816 704
rect 12256 756 12312 758
rect 12256 704 12258 756
rect 12258 704 12310 756
rect 12310 704 12312 756
rect 12256 702 12312 704
rect 14752 756 14808 758
rect 14752 704 14754 756
rect 14754 704 14806 756
rect 14806 704 14808 756
rect 14752 702 14808 704
rect 17248 756 17304 758
rect 17248 704 17250 756
rect 17250 704 17302 756
rect 17302 704 17304 756
rect 17248 702 17304 704
rect 19744 756 19800 758
rect 19744 704 19746 756
rect 19746 704 19798 756
rect 19798 704 19800 756
rect 19744 702 19800 704
rect 2272 434 2328 436
rect 2272 382 2274 434
rect 2274 382 2326 434
rect 2326 382 2328 434
rect 2272 380 2328 382
rect 4768 434 4824 436
rect 4768 382 4770 434
rect 4770 382 4822 434
rect 4822 382 4824 434
rect 4768 380 4824 382
rect 7264 434 7320 436
rect 7264 382 7266 434
rect 7266 382 7318 434
rect 7318 382 7320 434
rect 7264 380 7320 382
rect 9760 434 9816 436
rect 9760 382 9762 434
rect 9762 382 9814 434
rect 9814 382 9816 434
rect 9760 380 9816 382
rect 12256 434 12312 436
rect 12256 382 12258 434
rect 12258 382 12310 434
rect 12310 382 12312 434
rect 12256 380 12312 382
rect 14752 434 14808 436
rect 14752 382 14754 434
rect 14754 382 14806 434
rect 14806 382 14808 434
rect 14752 380 14808 382
rect 17248 434 17304 436
rect 17248 382 17250 434
rect 17250 382 17302 434
rect 17302 382 17304 434
rect 17248 380 17304 382
rect 19744 434 19800 436
rect 19744 382 19746 434
rect 19746 382 19798 434
rect 19798 382 19800 434
rect 19744 380 19800 382
<< metal3 >>
rect 2009 2524 2075 2527
rect 4505 2524 4571 2527
rect 7001 2524 7067 2527
rect 9497 2524 9563 2527
rect 11993 2524 12059 2527
rect 14489 2524 14555 2527
rect 16985 2524 17051 2527
rect 19481 2524 19547 2527
rect 0 2522 19891 2524
rect 0 2466 2014 2522
rect 2070 2466 4510 2522
rect 4566 2466 7006 2522
rect 7062 2466 9502 2522
rect 9558 2466 11998 2522
rect 12054 2466 14494 2522
rect 14550 2466 16990 2522
rect 17046 2466 19486 2522
rect 19542 2466 19891 2522
rect 0 2464 19891 2466
rect 2009 2461 2075 2464
rect 4505 2461 4571 2464
rect 7001 2461 7067 2464
rect 9497 2461 9563 2464
rect 11993 2461 12059 2464
rect 14489 2461 14555 2464
rect 16985 2461 17051 2464
rect 19481 2461 19547 2464
rect 33 2370 19924 2375
rect 33 2314 2342 2370
rect 2398 2314 4838 2370
rect 4894 2314 7334 2370
rect 7390 2314 9830 2370
rect 9886 2314 12326 2370
rect 12382 2314 14822 2370
rect 14878 2314 17318 2370
rect 17374 2314 19814 2370
rect 19870 2314 19924 2370
rect 33 2309 19924 2314
rect 33 1596 19924 1601
rect 33 1540 2260 1596
rect 2316 1540 4756 1596
rect 4812 1540 7252 1596
rect 7308 1540 9748 1596
rect 9804 1540 12244 1596
rect 12300 1540 14740 1596
rect 14796 1540 17236 1596
rect 17292 1540 19732 1596
rect 19788 1540 19924 1596
rect 33 1535 19924 1540
rect 33 758 19924 763
rect 33 702 2272 758
rect 2328 702 4768 758
rect 4824 702 7264 758
rect 7320 702 9760 758
rect 9816 702 12256 758
rect 12312 702 14752 758
rect 14808 702 17248 758
rect 17304 702 19744 758
rect 19800 702 19924 758
rect 33 697 19924 702
rect 33 436 19924 441
rect 33 380 2272 436
rect 2328 380 4768 436
rect 4824 380 7264 436
rect 7320 380 9760 436
rect 9816 380 12256 436
rect 12312 380 14752 436
rect 14808 380 17248 436
rect 17304 380 19744 436
rect 19800 380 19924 436
rect 33 375 19924 380
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1483185662
transform 1 0 19391 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1483185662
transform 1 0 16895 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1483185662
transform 1 0 14399 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1483185662
transform 1 0 11903 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1483185662
transform 1 0 9407 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1483185662
transform 1 0 6911 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1483185662
transform 1 0 4415 0 1 0
box -541 0 937 2556
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1483185662
transform 1 0 1919 0 1 0
box -541 0 937 2556
<< labels >>
rlabel metal1 s 2115 1430 2149 2556 4 bl_0
port 3 nsew
rlabel metal1 s 2191 1442 2219 2556 4 br_0
port 5 nsew
rlabel metal1 s 2023 0 2069 150 4 data_0
port 7 nsew
rlabel metal1 s 4611 1430 4645 2556 4 bl_1
port 9 nsew
rlabel metal1 s 4687 1442 4715 2556 4 br_1
port 11 nsew
rlabel metal1 s 4519 0 4565 150 4 data_1
port 13 nsew
rlabel metal1 s 7107 1430 7141 2556 4 bl_2
port 15 nsew
rlabel metal1 s 7183 1442 7211 2556 4 br_2
port 17 nsew
rlabel metal1 s 7015 0 7061 150 4 data_2
port 19 nsew
rlabel metal1 s 9603 1430 9637 2556 4 bl_3
port 21 nsew
rlabel metal1 s 9679 1442 9707 2556 4 br_3
port 23 nsew
rlabel metal1 s 9511 0 9557 150 4 data_3
port 25 nsew
rlabel metal1 s 12099 1430 12133 2556 4 bl_4
port 27 nsew
rlabel metal1 s 12175 1442 12203 2556 4 br_4
port 29 nsew
rlabel metal1 s 12007 0 12053 150 4 data_4
port 31 nsew
rlabel metal1 s 14595 1430 14629 2556 4 bl_5
port 33 nsew
rlabel metal1 s 14671 1442 14699 2556 4 br_5
port 35 nsew
rlabel metal1 s 14503 0 14549 150 4 data_5
port 37 nsew
rlabel metal1 s 17091 1430 17125 2556 4 bl_6
port 39 nsew
rlabel metal1 s 17167 1442 17195 2556 4 br_6
port 41 nsew
rlabel metal1 s 16999 0 17045 150 4 data_6
port 43 nsew
rlabel metal1 s 19587 1430 19621 2556 4 bl_7
port 45 nsew
rlabel metal1 s 19663 1442 19691 2556 4 br_7
port 47 nsew
rlabel metal1 s 19495 0 19541 150 4 data_7
port 49 nsew
rlabel metal3 s 33 1535 19924 1601 4 vdd
port 51 nsew
rlabel metal3 s 33 697 19924 763 4 vdd
port 51 nsew
rlabel metal3 s 33 375 19924 441 4 gnd
port 53 nsew
rlabel metal3 s 33 2309 19924 2375 4 gnd
port 53 nsew
rlabel metal3 s 0 2464 19891 2524 4 en
port 55 nsew
<< properties >>
string FIXED_BBOX 0 0 19891 2556
<< end >>
