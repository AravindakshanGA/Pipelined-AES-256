magic
tech sky130A
magscale 1 2
timestamp 1543373569
<< checkpaint >>
rect -1216 -1260 2020 1750
<< nwell >>
rect 428 0 760 490
<< pwell >>
rect 147 271 249 462
rect 136 69 260 271
<< scnmos >>
rect 162 155 234 185
<< scpmos >>
rect 482 155 706 185
<< ndiff >>
rect 162 237 234 245
rect 162 203 181 237
rect 215 203 234 237
rect 162 185 234 203
rect 162 137 234 155
rect 162 103 181 137
rect 215 103 234 137
rect 162 95 234 103
<< pdiff >>
rect 482 237 706 245
rect 482 203 577 237
rect 611 203 706 237
rect 482 185 706 203
rect 482 137 706 155
rect 482 103 577 137
rect 611 103 706 137
rect 482 95 706 103
<< ndiffc >>
rect 181 203 215 237
rect 181 103 215 137
<< pdiffc >>
rect 577 203 611 237
rect 577 103 611 137
<< psubdiff >>
rect 173 412 223 436
rect 173 378 181 412
rect 215 378 223 412
rect 173 354 223 378
<< nsubdiff >>
rect 569 412 619 436
rect 569 378 577 412
rect 611 378 619 412
rect 569 354 619 378
<< psubdiffcont >>
rect 181 378 215 412
<< nsubdiffcont >>
rect 577 378 611 412
<< poly >>
rect 44 187 110 203
rect 44 153 60 187
rect 94 185 110 187
rect 94 155 162 185
rect 234 155 482 185
rect 706 155 732 185
rect 94 153 110 155
rect 44 137 110 153
<< polycont >>
rect 60 153 94 187
<< locali >>
rect 181 412 215 428
rect 181 362 215 378
rect 577 412 611 428
rect 577 362 611 378
rect 181 237 215 253
rect 577 237 611 253
rect 165 203 181 237
rect 215 203 231 237
rect 561 203 577 237
rect 611 203 627 237
rect 60 187 94 203
rect 181 187 215 203
rect 577 187 611 203
rect 60 137 94 153
rect 165 103 181 137
rect 215 103 577 137
rect 611 103 742 137
<< viali >>
rect 181 378 215 412
rect 577 378 611 412
rect 181 203 215 237
rect 577 203 611 237
<< metal1 >>
rect 169 412 227 418
rect 169 378 181 412
rect 215 378 227 412
rect 169 372 227 378
rect 565 412 623 418
rect 565 378 577 412
rect 611 378 623 412
rect 565 372 623 378
rect 184 243 212 372
rect 580 243 608 372
rect 169 237 227 243
rect 169 203 181 237
rect 215 203 227 237
rect 169 197 227 203
rect 565 237 623 243
rect 565 203 577 237
rect 611 203 623 237
rect 565 197 623 203
rect 184 0 212 197
rect 580 0 608 197
<< labels >>
rlabel locali s 77 170 77 170 4 A
port 2 nsew
rlabel locali s 453 120 453 120 4 Z
port 3 nsew
rlabel metal1 s 184 0 212 395 4 gnd
port 5 nsew
rlabel metal1 s 580 0 608 395 4 vdd
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 742 41
<< end >>
