magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1309 3850 2731
<< locali >>
rect 1260 1432 1294 1447
rect 0 1431 2554 1432
rect 0 1397 1260 1431
rect 1294 1397 2554 1431
rect 0 1396 2554 1397
rect 1260 1381 1294 1396
rect 1260 18 1294 33
rect 0 17 2554 18
rect 0 -17 1260 17
rect 1294 -17 2554 17
rect 0 -18 2554 -17
rect 1260 -33 1294 -18
<< viali >>
rect 1260 1397 1294 1431
rect 1260 -17 1294 17
<< metal1 >>
rect 1245 1388 1251 1440
rect 1303 1388 1309 1440
rect 1245 -26 1251 26
rect 1303 -26 1309 26
<< via1 >>
rect 1251 1431 1303 1440
rect 1251 1397 1260 1431
rect 1260 1397 1294 1431
rect 1294 1397 1303 1431
rect 1251 1388 1303 1397
rect 1251 17 1303 26
rect 1251 -17 1260 17
rect 1260 -17 1294 17
rect 1294 -17 1303 17
rect 1251 -26 1303 -17
<< metal2 >>
rect 1249 1442 1305 1451
rect 137 538 203 590
rect 369 0 397 1414
rect 1249 1377 1305 1386
rect 1858 871 1886 899
rect 2364 489 2392 517
rect 1249 28 1305 37
rect 1249 -37 1305 -28
<< via2 >>
rect 1249 1440 1305 1442
rect 1249 1388 1251 1440
rect 1251 1388 1303 1440
rect 1303 1388 1305 1440
rect 1249 1386 1305 1388
rect 1249 26 1305 28
rect 1249 -26 1251 26
rect 1251 -26 1303 26
rect 1303 -26 1305 26
rect 1249 -28 1305 -26
<< metal3 >>
rect 1228 1442 1326 1463
rect 1228 1386 1249 1442
rect 1305 1386 1326 1442
rect 1228 1365 1326 1386
rect 1228 28 1326 49
rect 1228 -28 1249 28
rect 1305 -28 1326 28
rect 1228 -49 1326 -28
use subbyte2_dff_buf_0  subbyte2_dff_buf_0_0
timestamp 1543373571
transform 1 0 0 0 1 0
box -36 -43 2590 1471
<< labels >>
rlabel metal3 s 1228 1365 1326 1463 4 vdd
port 3 nsew
rlabel metal3 s 1228 -49 1326 49 4 gnd
port 5 nsew
rlabel metal2 s 137 538 203 590 4 din_0
port 7 nsew
rlabel metal2 s 2364 489 2392 517 4 dout_0
port 9 nsew
rlabel metal2 s 1858 871 1886 899 4 dout_bar_0
port 11 nsew
rlabel metal2 s 369 0 397 1414 4 clk
port 13 nsew
<< properties >>
string FIXED_BBOX 1244 -37 1310 0
<< end >>
