magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 1880 2731
<< nwell >>
rect -36 679 620 1471
<< pwell >>
rect 28 159 446 413
rect 28 25 550 159
<< scnmos >>
rect 114 51 144 387
rect 222 51 252 387
rect 330 51 360 387
<< scpmos >>
rect 114 1027 144 1363
rect 222 1027 252 1363
rect 330 1027 360 1363
<< ndiff >>
rect 54 236 114 387
rect 54 202 62 236
rect 96 202 114 236
rect 54 51 114 202
rect 144 236 222 387
rect 144 202 166 236
rect 200 202 222 236
rect 144 51 222 202
rect 252 236 330 387
rect 252 202 274 236
rect 308 202 330 236
rect 252 51 330 202
rect 360 236 420 387
rect 360 202 378 236
rect 412 202 420 236
rect 360 51 420 202
<< pdiff >>
rect 54 1212 114 1363
rect 54 1178 62 1212
rect 96 1178 114 1212
rect 54 1027 114 1178
rect 144 1212 222 1363
rect 144 1178 166 1212
rect 200 1178 222 1212
rect 144 1027 222 1178
rect 252 1212 330 1363
rect 252 1178 274 1212
rect 308 1178 330 1212
rect 252 1027 330 1178
rect 360 1212 420 1363
rect 360 1178 378 1212
rect 412 1178 420 1212
rect 360 1027 420 1178
<< ndiffc >>
rect 62 202 96 236
rect 166 202 200 236
rect 274 202 308 236
rect 378 202 412 236
<< pdiffc >>
rect 62 1178 96 1212
rect 166 1178 200 1212
rect 274 1178 308 1212
rect 378 1178 412 1212
<< psubdiff >>
rect 474 109 524 133
rect 474 75 482 109
rect 516 75 524 109
rect 474 51 524 75
<< nsubdiff >>
rect 474 1326 524 1350
rect 474 1292 482 1326
rect 516 1292 524 1326
rect 474 1268 524 1292
<< psubdiffcont >>
rect 482 75 516 109
<< nsubdiffcont >>
rect 482 1292 516 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 330 1363 360 1389
rect 114 1001 144 1027
rect 222 1001 252 1027
rect 330 1001 360 1027
rect 114 971 360 1001
rect 114 740 144 971
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 443 144 674
rect 114 413 360 443
rect 114 387 144 413
rect 222 387 252 413
rect 330 387 360 413
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 584 1431
rect 62 1212 96 1397
rect 62 1162 96 1178
rect 166 1212 200 1228
rect 166 1128 200 1178
rect 274 1212 308 1397
rect 482 1326 516 1397
rect 482 1276 516 1292
rect 274 1162 308 1178
rect 378 1212 412 1228
rect 378 1128 412 1178
rect 166 1094 412 1128
rect 64 724 98 740
rect 64 674 98 690
rect 272 724 306 1094
rect 272 690 323 724
rect 272 320 306 690
rect 166 286 412 320
rect 62 236 96 252
rect 62 17 96 202
rect 166 236 200 286
rect 166 186 200 202
rect 274 236 308 252
rect 274 17 308 202
rect 378 236 412 286
rect 378 186 412 202
rect 482 109 516 125
rect 482 17 516 75
rect 0 -17 584 17
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 306 707 306 707 4 Z
port 2 nsew
rlabel locali s 292 0 292 0 4 gnd
port 3 nsew
rlabel locali s 292 1414 292 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 584 1111
<< end >>
