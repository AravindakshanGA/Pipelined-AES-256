magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 2096 2731
<< nwell >>
rect -36 679 836 1471
<< pwell >>
rect 28 159 662 413
rect 28 25 766 159
<< scnmos >>
rect 114 51 144 387
rect 222 51 252 387
rect 330 51 360 387
rect 438 51 468 387
rect 546 51 576 387
<< scpmos >>
rect 114 963 144 1363
rect 222 963 252 1363
rect 330 963 360 1363
rect 438 963 468 1363
rect 546 963 576 1363
<< ndiff >>
rect 54 236 114 387
rect 54 202 62 236
rect 96 202 114 236
rect 54 51 114 202
rect 144 236 222 387
rect 144 202 166 236
rect 200 202 222 236
rect 144 51 222 202
rect 252 236 330 387
rect 252 202 274 236
rect 308 202 330 236
rect 252 51 330 202
rect 360 236 438 387
rect 360 202 382 236
rect 416 202 438 236
rect 360 51 438 202
rect 468 236 546 387
rect 468 202 490 236
rect 524 202 546 236
rect 468 51 546 202
rect 576 236 636 387
rect 576 202 594 236
rect 628 202 636 236
rect 576 51 636 202
<< pdiff >>
rect 54 1180 114 1363
rect 54 1146 62 1180
rect 96 1146 114 1180
rect 54 963 114 1146
rect 144 1180 222 1363
rect 144 1146 166 1180
rect 200 1146 222 1180
rect 144 963 222 1146
rect 252 1180 330 1363
rect 252 1146 274 1180
rect 308 1146 330 1180
rect 252 963 330 1146
rect 360 1180 438 1363
rect 360 1146 382 1180
rect 416 1146 438 1180
rect 360 963 438 1146
rect 468 1180 546 1363
rect 468 1146 490 1180
rect 524 1146 546 1180
rect 468 963 546 1146
rect 576 1180 636 1363
rect 576 1146 594 1180
rect 628 1146 636 1180
rect 576 963 636 1146
<< ndiffc >>
rect 62 202 96 236
rect 166 202 200 236
rect 274 202 308 236
rect 382 202 416 236
rect 490 202 524 236
rect 594 202 628 236
<< pdiffc >>
rect 62 1146 96 1180
rect 166 1146 200 1180
rect 274 1146 308 1180
rect 382 1146 416 1180
rect 490 1146 524 1180
rect 594 1146 628 1180
<< psubdiff >>
rect 690 109 740 133
rect 690 75 698 109
rect 732 75 740 109
rect 690 51 740 75
<< nsubdiff >>
rect 690 1326 740 1350
rect 690 1292 698 1326
rect 732 1292 740 1326
rect 690 1268 740 1292
<< psubdiffcont >>
rect 698 75 732 109
<< nsubdiffcont >>
rect 698 1292 732 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 330 1363 360 1389
rect 438 1363 468 1389
rect 546 1363 576 1389
rect 114 937 144 963
rect 222 937 252 963
rect 330 937 360 963
rect 438 937 468 963
rect 546 937 576 963
rect 114 907 576 937
rect 114 724 144 907
rect 48 708 144 724
rect 48 674 64 708
rect 98 674 144 708
rect 48 658 144 674
rect 114 443 144 658
rect 114 413 576 443
rect 114 387 144 413
rect 222 387 252 413
rect 330 387 360 413
rect 438 387 468 413
rect 546 387 576 413
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
<< polycont >>
rect 64 674 98 708
<< locali >>
rect 0 1397 800 1431
rect 62 1180 96 1397
rect 62 1130 96 1146
rect 166 1180 200 1196
rect 166 1096 200 1146
rect 274 1180 308 1397
rect 274 1130 308 1146
rect 382 1180 416 1196
rect 382 1096 416 1146
rect 490 1180 524 1397
rect 698 1326 732 1397
rect 698 1276 732 1292
rect 490 1130 524 1146
rect 594 1180 628 1196
rect 594 1096 628 1146
rect 166 1062 628 1096
rect 64 708 98 724
rect 64 658 98 674
rect 380 708 414 1062
rect 380 674 431 708
rect 380 320 414 674
rect 166 286 628 320
rect 62 236 96 252
rect 62 17 96 202
rect 166 236 200 286
rect 166 186 200 202
rect 274 236 308 252
rect 274 17 308 202
rect 382 236 416 286
rect 382 186 416 202
rect 490 236 524 252
rect 490 17 524 202
rect 594 236 628 286
rect 594 186 628 202
rect 698 109 732 125
rect 698 17 732 75
rect 0 -17 800 17
<< labels >>
rlabel locali s 81 691 81 691 4 A
port 1 nsew
rlabel locali s 414 691 414 691 4 Z
port 2 nsew
rlabel locali s 400 0 400 0 4 gnd
port 3 nsew
rlabel locali s 400 1414 400 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 800 1079
<< end >>
