magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1260 -1256 21531 3271
<< metal1 >>
rect 2045 1959 2075 2011
rect 2247 1959 2277 2011
rect 4541 1959 4571 2011
rect 4743 1959 4773 2011
rect 7037 1959 7067 2011
rect 7239 1959 7269 2011
rect 9533 1959 9563 2011
rect 9735 1959 9765 2011
rect 12029 1959 12059 2011
rect 12231 1959 12261 2011
rect 14525 1959 14555 2011
rect 14727 1959 14757 2011
rect 17021 1959 17051 2011
rect 17223 1959 17253 2011
rect 19517 1959 19547 2011
rect 19719 1959 19749 2011
rect 2154 1552 2160 1604
rect 2212 1552 2218 1604
rect 4650 1552 4656 1604
rect 4708 1552 4714 1604
rect 7146 1552 7152 1604
rect 7204 1552 7210 1604
rect 9642 1552 9648 1604
rect 9700 1552 9706 1604
rect 12138 1552 12144 1604
rect 12196 1552 12202 1604
rect 14634 1552 14640 1604
rect 14692 1552 14698 1604
rect 17130 1552 17136 1604
rect 17188 1552 17194 1604
rect 19626 1552 19632 1604
rect 19684 1552 19690 1604
rect 2143 1115 2149 1167
rect 2201 1115 2207 1167
rect 4639 1115 4645 1167
rect 4697 1115 4703 1167
rect 7135 1115 7141 1167
rect 7193 1115 7199 1167
rect 9631 1115 9637 1167
rect 9689 1115 9695 1167
rect 12127 1115 12133 1167
rect 12185 1115 12191 1167
rect 14623 1115 14629 1167
rect 14681 1115 14687 1167
rect 17119 1115 17125 1167
rect 17177 1115 17183 1167
rect 19615 1115 19621 1167
rect 19673 1115 19679 1167
rect 2264 784 2270 836
rect 2322 784 2328 836
rect 4760 784 4766 836
rect 4818 784 4824 836
rect 7256 784 7262 836
rect 7314 784 7320 836
rect 9752 784 9758 836
rect 9810 784 9816 836
rect 12248 784 12254 836
rect 12306 784 12312 836
rect 14744 784 14750 836
rect 14802 784 14808 836
rect 17240 784 17246 836
rect 17298 784 17304 836
rect 19736 784 19742 836
rect 19794 784 19800 836
rect 1987 291 1993 343
rect 2045 291 2051 343
rect 4483 291 4489 343
rect 4541 291 4547 343
rect 6979 291 6985 343
rect 7037 291 7043 343
rect 9475 291 9481 343
rect 9533 291 9539 343
rect 11971 291 11977 343
rect 12029 291 12035 343
rect 14467 291 14473 343
rect 14525 291 14531 343
rect 16963 291 16969 343
rect 17021 291 17027 343
rect 19459 291 19465 343
rect 19517 291 19523 343
rect 0 94 19891 122
rect 2142 4 2202 60
rect 4638 4 4698 60
rect 7134 4 7194 60
rect 9630 4 9690 60
rect 12126 4 12186 60
rect 14622 4 14682 60
rect 17118 4 17178 60
rect 19614 4 19674 60
<< via1 >>
rect 2160 1552 2212 1604
rect 4656 1552 4708 1604
rect 7152 1552 7204 1604
rect 9648 1552 9700 1604
rect 12144 1552 12196 1604
rect 14640 1552 14692 1604
rect 17136 1552 17188 1604
rect 19632 1552 19684 1604
rect 2149 1115 2201 1167
rect 4645 1115 4697 1167
rect 7141 1115 7193 1167
rect 9637 1115 9689 1167
rect 12133 1115 12185 1167
rect 14629 1115 14681 1167
rect 17125 1115 17177 1167
rect 19621 1115 19673 1167
rect 2270 784 2322 836
rect 4766 784 4818 836
rect 7262 784 7314 836
rect 9758 784 9810 836
rect 12254 784 12306 836
rect 14750 784 14802 836
rect 17246 784 17298 836
rect 19742 784 19794 836
rect 1993 291 2045 343
rect 4489 291 4541 343
rect 6985 291 7037 343
rect 9481 291 9533 343
rect 11977 291 12029 343
rect 14473 291 14525 343
rect 16969 291 17021 343
rect 19465 291 19517 343
<< metal2 >>
rect 2158 1606 2214 1615
rect 2158 1541 2214 1550
rect 4654 1606 4710 1615
rect 4654 1541 4710 1550
rect 7150 1606 7206 1615
rect 7150 1541 7206 1550
rect 9646 1606 9702 1615
rect 9646 1541 9702 1550
rect 12142 1606 12198 1615
rect 12142 1541 12198 1550
rect 14638 1606 14694 1615
rect 14638 1541 14694 1550
rect 17134 1606 17190 1615
rect 17134 1541 17190 1550
rect 19630 1606 19686 1615
rect 19630 1541 19686 1550
rect 2147 1169 2203 1178
rect 2147 1104 2203 1113
rect 4643 1169 4699 1178
rect 4643 1104 4699 1113
rect 7139 1169 7195 1178
rect 7139 1104 7195 1113
rect 9635 1169 9691 1178
rect 9635 1104 9691 1113
rect 12131 1169 12187 1178
rect 12131 1104 12187 1113
rect 14627 1169 14683 1178
rect 14627 1104 14683 1113
rect 17123 1169 17179 1178
rect 17123 1104 17179 1113
rect 19619 1169 19675 1178
rect 19619 1104 19675 1113
rect 2268 837 2324 846
rect 2268 772 2324 781
rect 4764 837 4820 846
rect 4764 772 4820 781
rect 7260 837 7316 846
rect 7260 772 7316 781
rect 9756 837 9812 846
rect 9756 772 9812 781
rect 12252 837 12308 846
rect 12252 772 12308 781
rect 14748 837 14804 846
rect 14748 772 14804 781
rect 17244 837 17300 846
rect 17244 772 17300 781
rect 19740 837 19796 846
rect 19740 772 19796 781
rect 1991 345 2047 354
rect 1991 280 2047 289
rect 4487 345 4543 354
rect 4487 280 4543 289
rect 6983 345 7039 354
rect 6983 280 7039 289
rect 9479 345 9535 354
rect 9479 280 9535 289
rect 11975 345 12031 354
rect 11975 280 12031 289
rect 14471 345 14527 354
rect 14471 280 14527 289
rect 16967 345 17023 354
rect 16967 280 17023 289
rect 19463 345 19519 354
rect 19463 280 19519 289
<< via2 >>
rect 2158 1604 2214 1606
rect 2158 1552 2160 1604
rect 2160 1552 2212 1604
rect 2212 1552 2214 1604
rect 2158 1550 2214 1552
rect 4654 1604 4710 1606
rect 4654 1552 4656 1604
rect 4656 1552 4708 1604
rect 4708 1552 4710 1604
rect 4654 1550 4710 1552
rect 7150 1604 7206 1606
rect 7150 1552 7152 1604
rect 7152 1552 7204 1604
rect 7204 1552 7206 1604
rect 7150 1550 7206 1552
rect 9646 1604 9702 1606
rect 9646 1552 9648 1604
rect 9648 1552 9700 1604
rect 9700 1552 9702 1604
rect 9646 1550 9702 1552
rect 12142 1604 12198 1606
rect 12142 1552 12144 1604
rect 12144 1552 12196 1604
rect 12196 1552 12198 1604
rect 12142 1550 12198 1552
rect 14638 1604 14694 1606
rect 14638 1552 14640 1604
rect 14640 1552 14692 1604
rect 14692 1552 14694 1604
rect 14638 1550 14694 1552
rect 17134 1604 17190 1606
rect 17134 1552 17136 1604
rect 17136 1552 17188 1604
rect 17188 1552 17190 1604
rect 17134 1550 17190 1552
rect 19630 1604 19686 1606
rect 19630 1552 19632 1604
rect 19632 1552 19684 1604
rect 19684 1552 19686 1604
rect 19630 1550 19686 1552
rect 2147 1167 2203 1169
rect 2147 1115 2149 1167
rect 2149 1115 2201 1167
rect 2201 1115 2203 1167
rect 2147 1113 2203 1115
rect 4643 1167 4699 1169
rect 4643 1115 4645 1167
rect 4645 1115 4697 1167
rect 4697 1115 4699 1167
rect 4643 1113 4699 1115
rect 7139 1167 7195 1169
rect 7139 1115 7141 1167
rect 7141 1115 7193 1167
rect 7193 1115 7195 1167
rect 7139 1113 7195 1115
rect 9635 1167 9691 1169
rect 9635 1115 9637 1167
rect 9637 1115 9689 1167
rect 9689 1115 9691 1167
rect 9635 1113 9691 1115
rect 12131 1167 12187 1169
rect 12131 1115 12133 1167
rect 12133 1115 12185 1167
rect 12185 1115 12187 1167
rect 12131 1113 12187 1115
rect 14627 1167 14683 1169
rect 14627 1115 14629 1167
rect 14629 1115 14681 1167
rect 14681 1115 14683 1167
rect 14627 1113 14683 1115
rect 17123 1167 17179 1169
rect 17123 1115 17125 1167
rect 17125 1115 17177 1167
rect 17177 1115 17179 1167
rect 17123 1113 17179 1115
rect 19619 1167 19675 1169
rect 19619 1115 19621 1167
rect 19621 1115 19673 1167
rect 19673 1115 19675 1167
rect 19619 1113 19675 1115
rect 2268 836 2324 837
rect 2268 784 2270 836
rect 2270 784 2322 836
rect 2322 784 2324 836
rect 2268 781 2324 784
rect 4764 836 4820 837
rect 4764 784 4766 836
rect 4766 784 4818 836
rect 4818 784 4820 836
rect 4764 781 4820 784
rect 7260 836 7316 837
rect 7260 784 7262 836
rect 7262 784 7314 836
rect 7314 784 7316 836
rect 7260 781 7316 784
rect 9756 836 9812 837
rect 9756 784 9758 836
rect 9758 784 9810 836
rect 9810 784 9812 836
rect 9756 781 9812 784
rect 12252 836 12308 837
rect 12252 784 12254 836
rect 12254 784 12306 836
rect 12306 784 12308 836
rect 12252 781 12308 784
rect 14748 836 14804 837
rect 14748 784 14750 836
rect 14750 784 14802 836
rect 14802 784 14804 836
rect 14748 781 14804 784
rect 17244 836 17300 837
rect 17244 784 17246 836
rect 17246 784 17298 836
rect 17298 784 17300 836
rect 17244 781 17300 784
rect 19740 836 19796 837
rect 19740 784 19742 836
rect 19742 784 19794 836
rect 19794 784 19796 836
rect 19740 781 19796 784
rect 1991 343 2047 345
rect 1991 291 1993 343
rect 1993 291 2045 343
rect 2045 291 2047 343
rect 1991 289 2047 291
rect 4487 343 4543 345
rect 4487 291 4489 343
rect 4489 291 4541 343
rect 4541 291 4543 343
rect 4487 289 4543 291
rect 6983 343 7039 345
rect 6983 291 6985 343
rect 6985 291 7037 343
rect 7037 291 7039 343
rect 6983 289 7039 291
rect 9479 343 9535 345
rect 9479 291 9481 343
rect 9481 291 9533 343
rect 9533 291 9535 343
rect 9479 289 9535 291
rect 11975 343 12031 345
rect 11975 291 11977 343
rect 11977 291 12029 343
rect 12029 291 12031 343
rect 11975 289 12031 291
rect 14471 343 14527 345
rect 14471 291 14473 343
rect 14473 291 14525 343
rect 14525 291 14527 343
rect 14471 289 14527 291
rect 16967 343 17023 345
rect 16967 291 16969 343
rect 16969 291 17021 343
rect 17021 291 17023 343
rect 16967 289 17023 291
rect 19463 343 19519 345
rect 19463 291 19465 343
rect 19465 291 19517 343
rect 19517 291 19519 343
rect 19463 289 19519 291
<< metal3 >>
rect 33 1606 19924 1611
rect 33 1550 2158 1606
rect 2214 1550 4654 1606
rect 4710 1550 7150 1606
rect 7206 1550 9646 1606
rect 9702 1550 12142 1606
rect 12198 1550 14638 1606
rect 14694 1550 17134 1606
rect 17190 1550 19630 1606
rect 19686 1550 19924 1606
rect 33 1545 19924 1550
rect 33 1169 19924 1174
rect 33 1113 2147 1169
rect 2203 1113 4643 1169
rect 4699 1113 7139 1169
rect 7195 1113 9635 1169
rect 9691 1113 12131 1169
rect 12187 1113 14627 1169
rect 14683 1113 17123 1169
rect 17179 1113 19619 1169
rect 19675 1113 19924 1169
rect 33 1108 19924 1113
rect 33 837 19924 842
rect 33 781 2268 837
rect 2324 781 4764 837
rect 4820 781 7260 837
rect 7316 781 9756 837
rect 9812 781 12252 837
rect 12308 781 14748 837
rect 14804 781 17244 837
rect 17300 781 19740 837
rect 19796 781 19924 837
rect 33 776 19924 781
rect 33 345 19924 350
rect 33 289 1991 345
rect 2047 289 4487 345
rect 4543 289 6983 345
rect 7039 289 9479 345
rect 9535 289 11975 345
rect 12031 289 14471 345
rect 14527 289 16967 345
rect 17023 289 19463 345
rect 19519 289 19924 345
rect 33 284 19924 289
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1480678001
transform 1 0 19391 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1480678001
transform 1 0 16895 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1480678001
transform 1 0 14399 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1480678001
transform 1 0 11903 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1480678001
transform 1 0 9407 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1480678001
transform 1 0 6911 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1480678001
transform 1 0 4415 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1480678001
transform 1 0 1919 0 1 0
box -376 4 880 2011
<< labels >>
rlabel metal1 s 2142 4 2202 60 4 data_0
port 3 nsew
rlabel metal1 s 2045 1959 2075 2011 4 bl_0
port 5 nsew
rlabel metal1 s 2247 1959 2277 2011 4 br_0
port 7 nsew
rlabel metal1 s 4638 4 4698 60 4 data_1
port 9 nsew
rlabel metal1 s 4541 1959 4571 2011 4 bl_1
port 11 nsew
rlabel metal1 s 4743 1959 4773 2011 4 br_1
port 13 nsew
rlabel metal1 s 7134 4 7194 60 4 data_2
port 15 nsew
rlabel metal1 s 7037 1959 7067 2011 4 bl_2
port 17 nsew
rlabel metal1 s 7239 1959 7269 2011 4 br_2
port 19 nsew
rlabel metal1 s 9630 4 9690 60 4 data_3
port 21 nsew
rlabel metal1 s 9533 1959 9563 2011 4 bl_3
port 23 nsew
rlabel metal1 s 9735 1959 9765 2011 4 br_3
port 25 nsew
rlabel metal1 s 12126 4 12186 60 4 data_4
port 27 nsew
rlabel metal1 s 12029 1959 12059 2011 4 bl_4
port 29 nsew
rlabel metal1 s 12231 1959 12261 2011 4 br_4
port 31 nsew
rlabel metal1 s 14622 4 14682 60 4 data_5
port 33 nsew
rlabel metal1 s 14525 1959 14555 2011 4 bl_5
port 35 nsew
rlabel metal1 s 14727 1959 14757 2011 4 br_5
port 37 nsew
rlabel metal1 s 17118 4 17178 60 4 data_6
port 39 nsew
rlabel metal1 s 17021 1959 17051 2011 4 bl_6
port 41 nsew
rlabel metal1 s 17223 1959 17253 2011 4 br_6
port 43 nsew
rlabel metal1 s 19614 4 19674 60 4 data_7
port 45 nsew
rlabel metal1 s 19517 1959 19547 2011 4 bl_7
port 47 nsew
rlabel metal1 s 19719 1959 19749 2011 4 br_7
port 49 nsew
rlabel metal1 s 0 94 19891 122 4 en
port 51 nsew
rlabel metal3 s 33 284 19924 350 4 vdd
port 53 nsew
rlabel metal3 s 33 1108 19924 1174 4 vdd
port 53 nsew
rlabel metal3 s 33 776 19924 842 4 gnd
port 55 nsew
rlabel metal3 s 33 1545 19924 1611 4 gnd
port 55 nsew
<< properties >>
string FIXED_BBOX 0 0 19891 2011
<< end >>
