magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 1772 2731
<< nwell >>
rect -36 679 512 1471
<< pwell >>
rect 28 159 338 225
rect 28 25 442 159
<< scnmos >>
rect 114 51 144 199
rect 222 51 252 199
<< scpmos >>
rect 114 1111 144 1363
rect 222 1111 252 1363
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 142 222 199
rect 144 108 166 142
rect 200 108 222 142
rect 144 51 222 108
rect 252 142 312 199
rect 252 108 270 142
rect 304 108 312 142
rect 252 51 312 108
<< pdiff >>
rect 54 1254 114 1363
rect 54 1220 62 1254
rect 96 1220 114 1254
rect 54 1111 114 1220
rect 144 1254 222 1363
rect 144 1220 166 1254
rect 200 1220 222 1254
rect 144 1111 222 1220
rect 252 1254 312 1363
rect 252 1220 270 1254
rect 304 1220 312 1254
rect 252 1111 312 1220
<< ndiffc >>
rect 62 108 96 142
rect 166 108 200 142
rect 270 108 304 142
<< pdiffc >>
rect 62 1220 96 1254
rect 166 1220 200 1254
rect 270 1220 304 1254
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 1326 416 1350
rect 366 1292 374 1326
rect 408 1292 416 1326
rect 366 1268 416 1292
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 1292 408 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 114 1085 144 1111
rect 222 1085 252 1111
rect 114 1055 252 1085
rect 114 714 144 1055
rect 48 698 144 714
rect 48 664 64 698
rect 98 664 144 698
rect 48 648 144 664
rect 114 255 144 648
rect 114 225 252 255
rect 114 199 144 225
rect 222 199 252 225
rect 114 25 144 51
rect 222 25 252 51
<< polycont >>
rect 64 664 98 698
<< locali >>
rect 0 1397 476 1431
rect 62 1254 96 1397
rect 62 1204 96 1220
rect 166 1254 200 1270
rect 64 698 98 714
rect 64 648 98 664
rect 166 698 200 1220
rect 270 1254 304 1397
rect 374 1326 408 1397
rect 374 1276 408 1292
rect 270 1204 304 1220
rect 166 664 217 698
rect 62 142 96 158
rect 62 17 96 108
rect 166 142 200 664
rect 166 92 200 108
rect 270 142 304 158
rect 270 17 304 108
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
<< labels >>
rlabel locali s 81 681 81 681 4 A
port 1 nsew
rlabel locali s 200 681 200 681 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 1414 238 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1153
<< end >>
