magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 1774 2731
<< nwell >>
rect -36 679 514 1471
<< pwell >>
rect 28 25 430 225
<< scnmos >>
rect 114 51 144 199
rect 214 51 244 199
rect 314 51 344 199
<< scpmos >>
rect 114 1139 144 1363
rect 214 1139 244 1363
rect 314 1139 344 1363
<< ndiff >>
rect 54 142 114 199
rect 54 108 62 142
rect 96 108 114 142
rect 54 51 114 108
rect 144 51 214 199
rect 244 51 314 199
rect 344 142 404 199
rect 344 108 362 142
rect 396 108 404 142
rect 344 51 404 108
<< pdiff >>
rect 54 1268 114 1363
rect 54 1234 62 1268
rect 96 1234 114 1268
rect 54 1139 114 1234
rect 144 1268 214 1363
rect 144 1234 162 1268
rect 196 1234 214 1268
rect 144 1139 214 1234
rect 244 1268 314 1363
rect 244 1234 262 1268
rect 296 1234 314 1268
rect 244 1139 314 1234
rect 344 1268 404 1363
rect 344 1234 362 1268
rect 396 1234 404 1268
rect 344 1139 404 1234
<< ndiffc >>
rect 62 108 96 142
rect 362 108 396 142
<< pdiffc >>
rect 62 1234 96 1268
rect 162 1234 196 1268
rect 262 1234 296 1268
rect 362 1234 396 1268
<< poly >>
rect 114 1363 144 1389
rect 214 1363 244 1389
rect 314 1363 344 1389
rect 114 303 144 1139
rect 214 427 244 1139
rect 314 551 344 1139
rect 314 535 395 551
rect 314 501 345 535
rect 379 501 395 535
rect 314 485 395 501
rect 196 411 262 427
rect 196 377 212 411
rect 246 377 262 411
rect 196 361 262 377
rect 63 287 144 303
rect 63 253 79 287
rect 113 253 144 287
rect 63 237 144 253
rect 114 199 144 237
rect 214 199 244 361
rect 314 199 344 485
rect 114 25 144 51
rect 214 25 244 51
rect 314 25 344 51
<< polycont >>
rect 345 501 379 535
rect 212 377 246 411
rect 79 253 113 287
<< locali >>
rect 0 1397 478 1431
rect 62 1268 96 1397
rect 62 1218 96 1234
rect 162 1268 196 1284
rect 162 1184 196 1234
rect 262 1268 296 1397
rect 262 1218 296 1234
rect 362 1268 396 1284
rect 362 1184 396 1234
rect 162 1150 464 1184
rect 345 535 379 551
rect 345 485 379 501
rect 212 411 246 427
rect 212 361 246 377
rect 79 287 113 303
rect 79 237 113 253
rect 430 158 464 1150
rect 62 142 96 158
rect 62 17 96 108
rect 362 142 464 158
rect 396 108 464 142
rect 362 92 464 108
rect 0 -17 478 17
<< labels >>
rlabel locali s 96 270 96 270 4 A
port 1 nsew
rlabel locali s 229 394 229 394 4 B
port 2 nsew
rlabel locali s 362 518 362 518 4 C
port 3 nsew
rlabel locali s 447 1167 447 1167 4 Z
port 4 nsew
rlabel locali s 239 0 239 0 4 gnd
port 5 nsew
rlabel locali s 239 1414 239 1414 4 vdd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 478 1167
<< end >>
