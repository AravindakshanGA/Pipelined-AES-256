magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 2852 2731
<< nwell >>
rect -36 679 1592 1471
<< pwell >>
rect 28 159 1418 477
rect 28 25 1522 159
<< scnmos >>
rect 114 51 144 451
rect 222 51 252 451
rect 330 51 360 451
rect 438 51 468 451
rect 546 51 576 451
rect 654 51 684 451
rect 762 51 792 451
rect 870 51 900 451
rect 978 51 1008 451
rect 1086 51 1116 451
rect 1194 51 1224 451
rect 1302 51 1332 451
<< scpmos >>
rect 114 963 144 1363
rect 222 963 252 1363
rect 330 963 360 1363
rect 438 963 468 1363
rect 546 963 576 1363
rect 654 963 684 1363
rect 762 963 792 1363
rect 870 963 900 1363
rect 978 963 1008 1363
rect 1086 963 1116 1363
rect 1194 963 1224 1363
rect 1302 963 1332 1363
<< ndiff >>
rect 54 268 114 451
rect 54 234 62 268
rect 96 234 114 268
rect 54 51 114 234
rect 144 268 222 451
rect 144 234 166 268
rect 200 234 222 268
rect 144 51 222 234
rect 252 268 330 451
rect 252 234 274 268
rect 308 234 330 268
rect 252 51 330 234
rect 360 268 438 451
rect 360 234 382 268
rect 416 234 438 268
rect 360 51 438 234
rect 468 268 546 451
rect 468 234 490 268
rect 524 234 546 268
rect 468 51 546 234
rect 576 268 654 451
rect 576 234 598 268
rect 632 234 654 268
rect 576 51 654 234
rect 684 268 762 451
rect 684 234 706 268
rect 740 234 762 268
rect 684 51 762 234
rect 792 268 870 451
rect 792 234 814 268
rect 848 234 870 268
rect 792 51 870 234
rect 900 268 978 451
rect 900 234 922 268
rect 956 234 978 268
rect 900 51 978 234
rect 1008 268 1086 451
rect 1008 234 1030 268
rect 1064 234 1086 268
rect 1008 51 1086 234
rect 1116 268 1194 451
rect 1116 234 1138 268
rect 1172 234 1194 268
rect 1116 51 1194 234
rect 1224 268 1302 451
rect 1224 234 1246 268
rect 1280 234 1302 268
rect 1224 51 1302 234
rect 1332 268 1392 451
rect 1332 234 1350 268
rect 1384 234 1392 268
rect 1332 51 1392 234
<< pdiff >>
rect 54 1180 114 1363
rect 54 1146 62 1180
rect 96 1146 114 1180
rect 54 963 114 1146
rect 144 1180 222 1363
rect 144 1146 166 1180
rect 200 1146 222 1180
rect 144 963 222 1146
rect 252 1180 330 1363
rect 252 1146 274 1180
rect 308 1146 330 1180
rect 252 963 330 1146
rect 360 1180 438 1363
rect 360 1146 382 1180
rect 416 1146 438 1180
rect 360 963 438 1146
rect 468 1180 546 1363
rect 468 1146 490 1180
rect 524 1146 546 1180
rect 468 963 546 1146
rect 576 1180 654 1363
rect 576 1146 598 1180
rect 632 1146 654 1180
rect 576 963 654 1146
rect 684 1180 762 1363
rect 684 1146 706 1180
rect 740 1146 762 1180
rect 684 963 762 1146
rect 792 1180 870 1363
rect 792 1146 814 1180
rect 848 1146 870 1180
rect 792 963 870 1146
rect 900 1180 978 1363
rect 900 1146 922 1180
rect 956 1146 978 1180
rect 900 963 978 1146
rect 1008 1180 1086 1363
rect 1008 1146 1030 1180
rect 1064 1146 1086 1180
rect 1008 963 1086 1146
rect 1116 1180 1194 1363
rect 1116 1146 1138 1180
rect 1172 1146 1194 1180
rect 1116 963 1194 1146
rect 1224 1180 1302 1363
rect 1224 1146 1246 1180
rect 1280 1146 1302 1180
rect 1224 963 1302 1146
rect 1332 1180 1392 1363
rect 1332 1146 1350 1180
rect 1384 1146 1392 1180
rect 1332 963 1392 1146
<< ndiffc >>
rect 62 234 96 268
rect 166 234 200 268
rect 274 234 308 268
rect 382 234 416 268
rect 490 234 524 268
rect 598 234 632 268
rect 706 234 740 268
rect 814 234 848 268
rect 922 234 956 268
rect 1030 234 1064 268
rect 1138 234 1172 268
rect 1246 234 1280 268
rect 1350 234 1384 268
<< pdiffc >>
rect 62 1146 96 1180
rect 166 1146 200 1180
rect 274 1146 308 1180
rect 382 1146 416 1180
rect 490 1146 524 1180
rect 598 1146 632 1180
rect 706 1146 740 1180
rect 814 1146 848 1180
rect 922 1146 956 1180
rect 1030 1146 1064 1180
rect 1138 1146 1172 1180
rect 1246 1146 1280 1180
rect 1350 1146 1384 1180
<< psubdiff >>
rect 1446 109 1496 133
rect 1446 75 1454 109
rect 1488 75 1496 109
rect 1446 51 1496 75
<< nsubdiff >>
rect 1446 1326 1496 1350
rect 1446 1292 1454 1326
rect 1488 1292 1496 1326
rect 1446 1268 1496 1292
<< psubdiffcont >>
rect 1454 75 1488 109
<< nsubdiffcont >>
rect 1454 1292 1488 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 330 1363 360 1389
rect 438 1363 468 1389
rect 546 1363 576 1389
rect 654 1363 684 1389
rect 762 1363 792 1389
rect 870 1363 900 1389
rect 978 1363 1008 1389
rect 1086 1363 1116 1389
rect 1194 1363 1224 1389
rect 1302 1363 1332 1389
rect 114 937 144 963
rect 222 937 252 963
rect 330 937 360 963
rect 438 937 468 963
rect 546 937 576 963
rect 654 937 684 963
rect 762 937 792 963
rect 870 937 900 963
rect 978 937 1008 963
rect 1086 937 1116 963
rect 1194 937 1224 963
rect 1302 937 1332 963
rect 114 907 1332 937
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
rect 114 477 1332 507
rect 114 451 144 477
rect 222 451 252 477
rect 330 451 360 477
rect 438 451 468 477
rect 546 451 576 477
rect 654 451 684 477
rect 762 451 792 477
rect 870 451 900 477
rect 978 451 1008 477
rect 1086 451 1116 477
rect 1194 451 1224 477
rect 1302 451 1332 477
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
rect 762 25 792 51
rect 870 25 900 51
rect 978 25 1008 51
rect 1086 25 1116 51
rect 1194 25 1224 51
rect 1302 25 1332 51
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1556 1431
rect 62 1180 96 1397
rect 62 1130 96 1146
rect 166 1180 200 1196
rect 166 1096 200 1146
rect 274 1180 308 1397
rect 274 1130 308 1146
rect 382 1180 416 1196
rect 382 1096 416 1146
rect 490 1180 524 1397
rect 490 1130 524 1146
rect 598 1180 632 1196
rect 598 1096 632 1146
rect 706 1180 740 1397
rect 706 1130 740 1146
rect 814 1180 848 1196
rect 814 1096 848 1146
rect 922 1180 956 1397
rect 922 1130 956 1146
rect 1030 1180 1064 1196
rect 1030 1096 1064 1146
rect 1138 1180 1172 1397
rect 1138 1130 1172 1146
rect 1246 1180 1280 1196
rect 1246 1096 1280 1146
rect 1350 1180 1384 1397
rect 1454 1326 1488 1397
rect 1454 1276 1488 1292
rect 1350 1130 1384 1146
rect 166 1062 1280 1096
rect 64 724 98 740
rect 64 674 98 690
rect 706 724 740 1062
rect 706 690 757 724
rect 706 352 740 690
rect 166 318 1280 352
rect 62 268 96 284
rect 62 17 96 234
rect 166 268 200 318
rect 166 218 200 234
rect 274 268 308 284
rect 274 17 308 234
rect 382 268 416 318
rect 382 218 416 234
rect 490 268 524 284
rect 490 17 524 234
rect 598 268 632 318
rect 598 218 632 234
rect 706 268 740 284
rect 706 17 740 234
rect 814 268 848 318
rect 814 218 848 234
rect 922 268 956 284
rect 922 17 956 234
rect 1030 268 1064 318
rect 1030 218 1064 234
rect 1138 268 1172 284
rect 1138 17 1172 234
rect 1246 268 1280 318
rect 1246 218 1280 234
rect 1350 268 1384 284
rect 1350 17 1384 234
rect 1454 109 1488 125
rect 1454 17 1488 75
rect 0 -17 1556 17
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 740 707 740 707 4 Z
port 2 nsew
rlabel locali s 778 0 778 0 4 gnd
port 3 nsew
rlabel locali s 778 1414 778 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1556 1079
<< end >>
