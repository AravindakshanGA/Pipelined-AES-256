magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -702 -1325 5088 26605
<< locali >>
rect 3782 25143 3816 25177
rect 574 25106 608 25122
rect 574 25056 608 25072
rect 558 24964 624 24998
rect 558 24772 624 24806
rect 574 24698 608 24714
rect 574 24648 608 24664
rect 3782 24593 3816 24627
rect 3782 24353 3816 24387
rect 574 24316 608 24332
rect 574 24266 608 24282
rect 558 24174 624 24208
rect 558 23982 624 24016
rect 574 23908 608 23924
rect 574 23858 608 23874
rect 3782 23803 3816 23837
rect 3782 23563 3816 23597
rect 574 23526 608 23542
rect 574 23476 608 23492
rect 558 23384 624 23418
rect 558 23192 624 23226
rect 574 23118 608 23134
rect 574 23068 608 23084
rect 3782 23013 3816 23047
rect 3782 22773 3816 22807
rect 574 22736 608 22752
rect 574 22686 608 22702
rect 558 22594 624 22628
rect 558 22402 624 22436
rect 574 22328 608 22344
rect 574 22278 608 22294
rect 3782 22223 3816 22257
rect 3782 21983 3816 22017
rect 574 21946 608 21962
rect 574 21896 608 21912
rect 558 21804 624 21838
rect 558 21612 624 21646
rect 574 21538 608 21554
rect 574 21488 608 21504
rect 3782 21433 3816 21467
rect 3782 21193 3816 21227
rect 574 21156 608 21172
rect 574 21106 608 21122
rect 558 21014 624 21048
rect 558 20822 624 20856
rect 574 20748 608 20764
rect 574 20698 608 20714
rect 3782 20643 3816 20677
rect 3782 20403 3816 20437
rect 574 20366 608 20382
rect 574 20316 608 20332
rect 558 20224 624 20258
rect 558 20032 624 20066
rect 574 19958 608 19974
rect 574 19908 608 19924
rect 3782 19853 3816 19887
rect 3782 19613 3816 19647
rect 574 19576 608 19592
rect 574 19526 608 19542
rect 558 19434 624 19468
rect 558 19242 624 19276
rect 574 19168 608 19184
rect 574 19118 608 19134
rect 3782 19063 3816 19097
rect 3782 18823 3816 18857
rect 574 18786 608 18802
rect 574 18736 608 18752
rect 558 18644 624 18678
rect 558 18452 624 18486
rect 574 18378 608 18394
rect 574 18328 608 18344
rect 3782 18273 3816 18307
rect 3782 18033 3816 18067
rect 574 17996 608 18012
rect 574 17946 608 17962
rect 558 17854 624 17888
rect 558 17662 624 17696
rect 574 17588 608 17604
rect 574 17538 608 17554
rect 3782 17483 3816 17517
rect 3782 17243 3816 17277
rect 574 17206 608 17222
rect 574 17156 608 17172
rect 558 17064 624 17098
rect 558 16872 624 16906
rect 574 16798 608 16814
rect 574 16748 608 16764
rect 3782 16693 3816 16727
rect 3782 16453 3816 16487
rect 574 16416 608 16432
rect 574 16366 608 16382
rect 558 16274 624 16308
rect 558 16082 624 16116
rect 574 16008 608 16024
rect 574 15958 608 15974
rect 3782 15903 3816 15937
rect 3782 15663 3816 15697
rect 574 15626 608 15642
rect 574 15576 608 15592
rect 558 15484 624 15518
rect 558 15292 624 15326
rect 574 15218 608 15234
rect 574 15168 608 15184
rect 3782 15113 3816 15147
rect 3782 14873 3816 14907
rect 574 14836 608 14852
rect 574 14786 608 14802
rect 558 14694 624 14728
rect 558 14502 624 14536
rect 574 14428 608 14444
rect 574 14378 608 14394
rect 3782 14323 3816 14357
rect 3782 14083 3816 14117
rect 574 14046 608 14062
rect 574 13996 608 14012
rect 558 13904 624 13938
rect 558 13712 624 13746
rect 574 13638 608 13654
rect 574 13588 608 13604
rect 3782 13533 3816 13567
rect 3782 13293 3816 13327
rect 574 13256 608 13272
rect 574 13206 608 13222
rect 558 13114 624 13148
rect 558 12922 624 12956
rect 574 12848 608 12864
rect 574 12798 608 12814
rect 3782 12743 3816 12777
rect 3782 12503 3816 12537
rect 574 12466 608 12482
rect 574 12416 608 12432
rect 558 12324 624 12358
rect 558 12132 624 12166
rect 574 12058 608 12074
rect 574 12008 608 12024
rect 3782 11953 3816 11987
rect 3782 11713 3816 11747
rect 574 11676 608 11692
rect 574 11626 608 11642
rect 558 11534 624 11568
rect 558 11342 624 11376
rect 574 11268 608 11284
rect 574 11218 608 11234
rect 3782 11163 3816 11197
rect 3782 10923 3816 10957
rect 574 10886 608 10902
rect 574 10836 608 10852
rect 558 10744 624 10778
rect 558 10552 624 10586
rect 574 10478 608 10494
rect 574 10428 608 10444
rect 3782 10373 3816 10407
rect 3782 10133 3816 10167
rect 574 10096 608 10112
rect 574 10046 608 10062
rect 558 9954 624 9988
rect 558 9762 624 9796
rect 574 9688 608 9704
rect 574 9638 608 9654
rect 3782 9583 3816 9617
rect 3782 9343 3816 9377
rect 574 9306 608 9322
rect 574 9256 608 9272
rect 558 9164 624 9198
rect 558 8972 624 9006
rect 574 8898 608 8914
rect 574 8848 608 8864
rect 3782 8793 3816 8827
rect 3782 8553 3816 8587
rect 574 8516 608 8532
rect 574 8466 608 8482
rect 558 8374 624 8408
rect 558 8182 624 8216
rect 574 8108 608 8124
rect 574 8058 608 8074
rect 3782 8003 3816 8037
rect 3782 7763 3816 7797
rect 574 7726 608 7742
rect 574 7676 608 7692
rect 558 7584 624 7618
rect 558 7392 624 7426
rect 574 7318 608 7334
rect 574 7268 608 7284
rect 3782 7213 3816 7247
rect 3782 6973 3816 7007
rect 574 6936 608 6952
rect 574 6886 608 6902
rect 558 6794 624 6828
rect 558 6602 624 6636
rect 574 6528 608 6544
rect 574 6478 608 6494
rect 3782 6423 3816 6457
rect 3782 6183 3816 6217
rect 574 6146 608 6162
rect 574 6096 608 6112
rect 558 6004 624 6038
rect 558 5812 624 5846
rect 574 5738 608 5754
rect 574 5688 608 5704
rect 3782 5633 3816 5667
rect 3782 5393 3816 5427
rect 574 5356 608 5372
rect 574 5306 608 5322
rect 558 5214 624 5248
rect 558 5022 624 5056
rect 574 4948 608 4964
rect 574 4898 608 4914
rect 3782 4843 3816 4877
rect 3782 4603 3816 4637
rect 574 4566 608 4582
rect 574 4516 608 4532
rect 558 4424 624 4458
rect 558 4232 624 4266
rect 574 4158 608 4174
rect 574 4108 608 4124
rect 3782 4053 3816 4087
rect 3782 3813 3816 3847
rect 574 3776 608 3792
rect 574 3726 608 3742
rect 558 3634 624 3668
rect 558 3442 624 3476
rect 574 3368 608 3384
rect 574 3318 608 3334
rect 3782 3263 3816 3297
rect 3782 3023 3816 3057
rect 574 2986 608 3002
rect 574 2936 608 2952
rect 558 2844 624 2878
rect 558 2652 624 2686
rect 574 2578 608 2594
rect 574 2528 608 2544
rect 3782 2473 3816 2507
rect 3782 2233 3816 2267
rect 574 2196 608 2212
rect 574 2146 608 2162
rect 558 2054 624 2088
rect 558 1862 624 1896
rect 574 1788 608 1804
rect 574 1738 608 1754
rect 3782 1683 3816 1717
rect 3782 1443 3816 1477
rect 574 1406 608 1422
rect 574 1356 608 1372
rect 558 1264 624 1298
rect 558 1072 624 1106
rect 574 998 608 1014
rect 574 948 608 964
rect 3782 893 3816 927
rect 3782 653 3816 687
rect 574 616 608 632
rect 574 566 608 582
rect 558 474 624 508
rect 558 282 624 316
rect 574 208 608 224
rect 574 158 608 174
rect 3782 103 3816 137
<< viali >>
rect 574 25072 608 25106
rect 574 24664 608 24698
rect 574 24282 608 24316
rect 574 23874 608 23908
rect 574 23492 608 23526
rect 574 23084 608 23118
rect 574 22702 608 22736
rect 574 22294 608 22328
rect 574 21912 608 21946
rect 574 21504 608 21538
rect 574 21122 608 21156
rect 574 20714 608 20748
rect 574 20332 608 20366
rect 574 19924 608 19958
rect 574 19542 608 19576
rect 574 19134 608 19168
rect 574 18752 608 18786
rect 574 18344 608 18378
rect 574 17962 608 17996
rect 574 17554 608 17588
rect 574 17172 608 17206
rect 574 16764 608 16798
rect 574 16382 608 16416
rect 574 15974 608 16008
rect 574 15592 608 15626
rect 574 15184 608 15218
rect 574 14802 608 14836
rect 574 14394 608 14428
rect 574 14012 608 14046
rect 574 13604 608 13638
rect 574 13222 608 13256
rect 574 12814 608 12848
rect 574 12432 608 12466
rect 574 12024 608 12058
rect 574 11642 608 11676
rect 574 11234 608 11268
rect 574 10852 608 10886
rect 574 10444 608 10478
rect 574 10062 608 10096
rect 574 9654 608 9688
rect 574 9272 608 9306
rect 574 8864 608 8898
rect 574 8482 608 8516
rect 574 8074 608 8108
rect 574 7692 608 7726
rect 574 7284 608 7318
rect 574 6902 608 6936
rect 574 6494 608 6528
rect 574 6112 608 6146
rect 574 5704 608 5738
rect 574 5322 608 5356
rect 574 4914 608 4948
rect 574 4532 608 4566
rect 574 4124 608 4158
rect 574 3742 608 3776
rect 574 3334 608 3368
rect 574 2952 608 2986
rect 574 2544 608 2578
rect 574 2162 608 2196
rect 574 1754 608 1788
rect 574 1372 608 1406
rect 574 964 608 998
rect 574 582 608 616
rect 574 174 608 208
<< metal1 >>
rect 559 25063 565 25115
rect 617 25063 623 25115
rect 726 25068 732 25120
rect 784 25068 790 25120
rect 1151 25069 1157 25121
rect 1209 25069 1215 25121
rect 1794 25056 1800 25108
rect 1852 25056 1858 25108
rect 3042 25056 3048 25108
rect 3100 25056 3106 25108
rect 559 24655 565 24707
rect 617 24655 623 24707
rect 726 24650 732 24702
rect 784 24650 790 24702
rect 1151 24649 1157 24701
rect 1209 24649 1215 24701
rect 1794 24662 1800 24714
rect 1852 24662 1858 24714
rect 3042 24662 3048 24714
rect 3100 24662 3106 24714
rect 559 24273 565 24325
rect 617 24273 623 24325
rect 726 24278 732 24330
rect 784 24278 790 24330
rect 1151 24279 1157 24331
rect 1209 24279 1215 24331
rect 1794 24266 1800 24318
rect 1852 24266 1858 24318
rect 3042 24266 3048 24318
rect 3100 24266 3106 24318
rect 559 23865 565 23917
rect 617 23865 623 23917
rect 726 23860 732 23912
rect 784 23860 790 23912
rect 1151 23859 1157 23911
rect 1209 23859 1215 23911
rect 1794 23872 1800 23924
rect 1852 23872 1858 23924
rect 3042 23872 3048 23924
rect 3100 23872 3106 23924
rect 559 23483 565 23535
rect 617 23483 623 23535
rect 726 23488 732 23540
rect 784 23488 790 23540
rect 1151 23489 1157 23541
rect 1209 23489 1215 23541
rect 1794 23476 1800 23528
rect 1852 23476 1858 23528
rect 3042 23476 3048 23528
rect 3100 23476 3106 23528
rect 559 23075 565 23127
rect 617 23075 623 23127
rect 726 23070 732 23122
rect 784 23070 790 23122
rect 1151 23069 1157 23121
rect 1209 23069 1215 23121
rect 1794 23082 1800 23134
rect 1852 23082 1858 23134
rect 3042 23082 3048 23134
rect 3100 23082 3106 23134
rect 559 22693 565 22745
rect 617 22693 623 22745
rect 726 22698 732 22750
rect 784 22698 790 22750
rect 1151 22699 1157 22751
rect 1209 22699 1215 22751
rect 1794 22686 1800 22738
rect 1852 22686 1858 22738
rect 3042 22686 3048 22738
rect 3100 22686 3106 22738
rect 559 22285 565 22337
rect 617 22285 623 22337
rect 726 22280 732 22332
rect 784 22280 790 22332
rect 1151 22279 1157 22331
rect 1209 22279 1215 22331
rect 1794 22292 1800 22344
rect 1852 22292 1858 22344
rect 3042 22292 3048 22344
rect 3100 22292 3106 22344
rect 559 21903 565 21955
rect 617 21903 623 21955
rect 726 21908 732 21960
rect 784 21908 790 21960
rect 1151 21909 1157 21961
rect 1209 21909 1215 21961
rect 1794 21896 1800 21948
rect 1852 21896 1858 21948
rect 3042 21896 3048 21948
rect 3100 21896 3106 21948
rect 559 21495 565 21547
rect 617 21495 623 21547
rect 726 21490 732 21542
rect 784 21490 790 21542
rect 1151 21489 1157 21541
rect 1209 21489 1215 21541
rect 1794 21502 1800 21554
rect 1852 21502 1858 21554
rect 3042 21502 3048 21554
rect 3100 21502 3106 21554
rect 559 21113 565 21165
rect 617 21113 623 21165
rect 726 21118 732 21170
rect 784 21118 790 21170
rect 1151 21119 1157 21171
rect 1209 21119 1215 21171
rect 1794 21106 1800 21158
rect 1852 21106 1858 21158
rect 3042 21106 3048 21158
rect 3100 21106 3106 21158
rect 559 20705 565 20757
rect 617 20705 623 20757
rect 726 20700 732 20752
rect 784 20700 790 20752
rect 1151 20699 1157 20751
rect 1209 20699 1215 20751
rect 1794 20712 1800 20764
rect 1852 20712 1858 20764
rect 3042 20712 3048 20764
rect 3100 20712 3106 20764
rect 559 20323 565 20375
rect 617 20323 623 20375
rect 726 20328 732 20380
rect 784 20328 790 20380
rect 1151 20329 1157 20381
rect 1209 20329 1215 20381
rect 1794 20316 1800 20368
rect 1852 20316 1858 20368
rect 3042 20316 3048 20368
rect 3100 20316 3106 20368
rect 559 19915 565 19967
rect 617 19915 623 19967
rect 726 19910 732 19962
rect 784 19910 790 19962
rect 1151 19909 1157 19961
rect 1209 19909 1215 19961
rect 1794 19922 1800 19974
rect 1852 19922 1858 19974
rect 3042 19922 3048 19974
rect 3100 19922 3106 19974
rect 559 19533 565 19585
rect 617 19533 623 19585
rect 726 19538 732 19590
rect 784 19538 790 19590
rect 1151 19539 1157 19591
rect 1209 19539 1215 19591
rect 1794 19526 1800 19578
rect 1852 19526 1858 19578
rect 3042 19526 3048 19578
rect 3100 19526 3106 19578
rect 559 19125 565 19177
rect 617 19125 623 19177
rect 726 19120 732 19172
rect 784 19120 790 19172
rect 1151 19119 1157 19171
rect 1209 19119 1215 19171
rect 1794 19132 1800 19184
rect 1852 19132 1858 19184
rect 3042 19132 3048 19184
rect 3100 19132 3106 19184
rect 559 18743 565 18795
rect 617 18743 623 18795
rect 726 18748 732 18800
rect 784 18748 790 18800
rect 1151 18749 1157 18801
rect 1209 18749 1215 18801
rect 1794 18736 1800 18788
rect 1852 18736 1858 18788
rect 3042 18736 3048 18788
rect 3100 18736 3106 18788
rect 559 18335 565 18387
rect 617 18335 623 18387
rect 726 18330 732 18382
rect 784 18330 790 18382
rect 1151 18329 1157 18381
rect 1209 18329 1215 18381
rect 1794 18342 1800 18394
rect 1852 18342 1858 18394
rect 3042 18342 3048 18394
rect 3100 18342 3106 18394
rect 559 17953 565 18005
rect 617 17953 623 18005
rect 726 17958 732 18010
rect 784 17958 790 18010
rect 1151 17959 1157 18011
rect 1209 17959 1215 18011
rect 1794 17946 1800 17998
rect 1852 17946 1858 17998
rect 3042 17946 3048 17998
rect 3100 17946 3106 17998
rect 559 17545 565 17597
rect 617 17545 623 17597
rect 726 17540 732 17592
rect 784 17540 790 17592
rect 1151 17539 1157 17591
rect 1209 17539 1215 17591
rect 1794 17552 1800 17604
rect 1852 17552 1858 17604
rect 3042 17552 3048 17604
rect 3100 17552 3106 17604
rect 559 17163 565 17215
rect 617 17163 623 17215
rect 726 17168 732 17220
rect 784 17168 790 17220
rect 1151 17169 1157 17221
rect 1209 17169 1215 17221
rect 1794 17156 1800 17208
rect 1852 17156 1858 17208
rect 3042 17156 3048 17208
rect 3100 17156 3106 17208
rect 559 16755 565 16807
rect 617 16755 623 16807
rect 726 16750 732 16802
rect 784 16750 790 16802
rect 1151 16749 1157 16801
rect 1209 16749 1215 16801
rect 1794 16762 1800 16814
rect 1852 16762 1858 16814
rect 3042 16762 3048 16814
rect 3100 16762 3106 16814
rect 559 16373 565 16425
rect 617 16373 623 16425
rect 726 16378 732 16430
rect 784 16378 790 16430
rect 1151 16379 1157 16431
rect 1209 16379 1215 16431
rect 1794 16366 1800 16418
rect 1852 16366 1858 16418
rect 3042 16366 3048 16418
rect 3100 16366 3106 16418
rect 559 15965 565 16017
rect 617 15965 623 16017
rect 726 15960 732 16012
rect 784 15960 790 16012
rect 1151 15959 1157 16011
rect 1209 15959 1215 16011
rect 1794 15972 1800 16024
rect 1852 15972 1858 16024
rect 3042 15972 3048 16024
rect 3100 15972 3106 16024
rect 559 15583 565 15635
rect 617 15583 623 15635
rect 726 15588 732 15640
rect 784 15588 790 15640
rect 1151 15589 1157 15641
rect 1209 15589 1215 15641
rect 1794 15576 1800 15628
rect 1852 15576 1858 15628
rect 3042 15576 3048 15628
rect 3100 15576 3106 15628
rect 559 15175 565 15227
rect 617 15175 623 15227
rect 726 15170 732 15222
rect 784 15170 790 15222
rect 1151 15169 1157 15221
rect 1209 15169 1215 15221
rect 1794 15182 1800 15234
rect 1852 15182 1858 15234
rect 3042 15182 3048 15234
rect 3100 15182 3106 15234
rect 559 14793 565 14845
rect 617 14793 623 14845
rect 726 14798 732 14850
rect 784 14798 790 14850
rect 1151 14799 1157 14851
rect 1209 14799 1215 14851
rect 1794 14786 1800 14838
rect 1852 14786 1858 14838
rect 3042 14786 3048 14838
rect 3100 14786 3106 14838
rect 559 14385 565 14437
rect 617 14385 623 14437
rect 726 14380 732 14432
rect 784 14380 790 14432
rect 1151 14379 1157 14431
rect 1209 14379 1215 14431
rect 1794 14392 1800 14444
rect 1852 14392 1858 14444
rect 3042 14392 3048 14444
rect 3100 14392 3106 14444
rect 559 14003 565 14055
rect 617 14003 623 14055
rect 726 14008 732 14060
rect 784 14008 790 14060
rect 1151 14009 1157 14061
rect 1209 14009 1215 14061
rect 1794 13996 1800 14048
rect 1852 13996 1858 14048
rect 3042 13996 3048 14048
rect 3100 13996 3106 14048
rect 559 13595 565 13647
rect 617 13595 623 13647
rect 726 13590 732 13642
rect 784 13590 790 13642
rect 1151 13589 1157 13641
rect 1209 13589 1215 13641
rect 1794 13602 1800 13654
rect 1852 13602 1858 13654
rect 3042 13602 3048 13654
rect 3100 13602 3106 13654
rect 559 13213 565 13265
rect 617 13213 623 13265
rect 726 13218 732 13270
rect 784 13218 790 13270
rect 1151 13219 1157 13271
rect 1209 13219 1215 13271
rect 1794 13206 1800 13258
rect 1852 13206 1858 13258
rect 3042 13206 3048 13258
rect 3100 13206 3106 13258
rect 559 12805 565 12857
rect 617 12805 623 12857
rect 726 12800 732 12852
rect 784 12800 790 12852
rect 1151 12799 1157 12851
rect 1209 12799 1215 12851
rect 1794 12812 1800 12864
rect 1852 12812 1858 12864
rect 3042 12812 3048 12864
rect 3100 12812 3106 12864
rect 559 12423 565 12475
rect 617 12423 623 12475
rect 726 12428 732 12480
rect 784 12428 790 12480
rect 1151 12429 1157 12481
rect 1209 12429 1215 12481
rect 1794 12416 1800 12468
rect 1852 12416 1858 12468
rect 3042 12416 3048 12468
rect 3100 12416 3106 12468
rect 559 12015 565 12067
rect 617 12015 623 12067
rect 726 12010 732 12062
rect 784 12010 790 12062
rect 1151 12009 1157 12061
rect 1209 12009 1215 12061
rect 1794 12022 1800 12074
rect 1852 12022 1858 12074
rect 3042 12022 3048 12074
rect 3100 12022 3106 12074
rect 559 11633 565 11685
rect 617 11633 623 11685
rect 726 11638 732 11690
rect 784 11638 790 11690
rect 1151 11639 1157 11691
rect 1209 11639 1215 11691
rect 1794 11626 1800 11678
rect 1852 11626 1858 11678
rect 3042 11626 3048 11678
rect 3100 11626 3106 11678
rect 559 11225 565 11277
rect 617 11225 623 11277
rect 726 11220 732 11272
rect 784 11220 790 11272
rect 1151 11219 1157 11271
rect 1209 11219 1215 11271
rect 1794 11232 1800 11284
rect 1852 11232 1858 11284
rect 3042 11232 3048 11284
rect 3100 11232 3106 11284
rect 559 10843 565 10895
rect 617 10843 623 10895
rect 726 10848 732 10900
rect 784 10848 790 10900
rect 1151 10849 1157 10901
rect 1209 10849 1215 10901
rect 1794 10836 1800 10888
rect 1852 10836 1858 10888
rect 3042 10836 3048 10888
rect 3100 10836 3106 10888
rect 559 10435 565 10487
rect 617 10435 623 10487
rect 726 10430 732 10482
rect 784 10430 790 10482
rect 1151 10429 1157 10481
rect 1209 10429 1215 10481
rect 1794 10442 1800 10494
rect 1852 10442 1858 10494
rect 3042 10442 3048 10494
rect 3100 10442 3106 10494
rect 559 10053 565 10105
rect 617 10053 623 10105
rect 726 10058 732 10110
rect 784 10058 790 10110
rect 1151 10059 1157 10111
rect 1209 10059 1215 10111
rect 1794 10046 1800 10098
rect 1852 10046 1858 10098
rect 3042 10046 3048 10098
rect 3100 10046 3106 10098
rect 559 9645 565 9697
rect 617 9645 623 9697
rect 726 9640 732 9692
rect 784 9640 790 9692
rect 1151 9639 1157 9691
rect 1209 9639 1215 9691
rect 1794 9652 1800 9704
rect 1852 9652 1858 9704
rect 3042 9652 3048 9704
rect 3100 9652 3106 9704
rect 559 9263 565 9315
rect 617 9263 623 9315
rect 726 9268 732 9320
rect 784 9268 790 9320
rect 1151 9269 1157 9321
rect 1209 9269 1215 9321
rect 1794 9256 1800 9308
rect 1852 9256 1858 9308
rect 3042 9256 3048 9308
rect 3100 9256 3106 9308
rect 559 8855 565 8907
rect 617 8855 623 8907
rect 726 8850 732 8902
rect 784 8850 790 8902
rect 1151 8849 1157 8901
rect 1209 8849 1215 8901
rect 1794 8862 1800 8914
rect 1852 8862 1858 8914
rect 3042 8862 3048 8914
rect 3100 8862 3106 8914
rect 559 8473 565 8525
rect 617 8473 623 8525
rect 726 8478 732 8530
rect 784 8478 790 8530
rect 1151 8479 1157 8531
rect 1209 8479 1215 8531
rect 1794 8466 1800 8518
rect 1852 8466 1858 8518
rect 3042 8466 3048 8518
rect 3100 8466 3106 8518
rect 559 8065 565 8117
rect 617 8065 623 8117
rect 726 8060 732 8112
rect 784 8060 790 8112
rect 1151 8059 1157 8111
rect 1209 8059 1215 8111
rect 1794 8072 1800 8124
rect 1852 8072 1858 8124
rect 3042 8072 3048 8124
rect 3100 8072 3106 8124
rect 559 7683 565 7735
rect 617 7683 623 7735
rect 726 7688 732 7740
rect 784 7688 790 7740
rect 1151 7689 1157 7741
rect 1209 7689 1215 7741
rect 1794 7676 1800 7728
rect 1852 7676 1858 7728
rect 3042 7676 3048 7728
rect 3100 7676 3106 7728
rect 559 7275 565 7327
rect 617 7275 623 7327
rect 726 7270 732 7322
rect 784 7270 790 7322
rect 1151 7269 1157 7321
rect 1209 7269 1215 7321
rect 1794 7282 1800 7334
rect 1852 7282 1858 7334
rect 3042 7282 3048 7334
rect 3100 7282 3106 7334
rect 559 6893 565 6945
rect 617 6893 623 6945
rect 726 6898 732 6950
rect 784 6898 790 6950
rect 1151 6899 1157 6951
rect 1209 6899 1215 6951
rect 1794 6886 1800 6938
rect 1852 6886 1858 6938
rect 3042 6886 3048 6938
rect 3100 6886 3106 6938
rect 559 6485 565 6537
rect 617 6485 623 6537
rect 726 6480 732 6532
rect 784 6480 790 6532
rect 1151 6479 1157 6531
rect 1209 6479 1215 6531
rect 1794 6492 1800 6544
rect 1852 6492 1858 6544
rect 3042 6492 3048 6544
rect 3100 6492 3106 6544
rect 559 6103 565 6155
rect 617 6103 623 6155
rect 726 6108 732 6160
rect 784 6108 790 6160
rect 1151 6109 1157 6161
rect 1209 6109 1215 6161
rect 1794 6096 1800 6148
rect 1852 6096 1858 6148
rect 3042 6096 3048 6148
rect 3100 6096 3106 6148
rect 559 5695 565 5747
rect 617 5695 623 5747
rect 726 5690 732 5742
rect 784 5690 790 5742
rect 1151 5689 1157 5741
rect 1209 5689 1215 5741
rect 1794 5702 1800 5754
rect 1852 5702 1858 5754
rect 3042 5702 3048 5754
rect 3100 5702 3106 5754
rect 559 5313 565 5365
rect 617 5313 623 5365
rect 726 5318 732 5370
rect 784 5318 790 5370
rect 1151 5319 1157 5371
rect 1209 5319 1215 5371
rect 1794 5306 1800 5358
rect 1852 5306 1858 5358
rect 3042 5306 3048 5358
rect 3100 5306 3106 5358
rect 559 4905 565 4957
rect 617 4905 623 4957
rect 726 4900 732 4952
rect 784 4900 790 4952
rect 1151 4899 1157 4951
rect 1209 4899 1215 4951
rect 1794 4912 1800 4964
rect 1852 4912 1858 4964
rect 3042 4912 3048 4964
rect 3100 4912 3106 4964
rect 559 4523 565 4575
rect 617 4523 623 4575
rect 726 4528 732 4580
rect 784 4528 790 4580
rect 1151 4529 1157 4581
rect 1209 4529 1215 4581
rect 1794 4516 1800 4568
rect 1852 4516 1858 4568
rect 3042 4516 3048 4568
rect 3100 4516 3106 4568
rect 559 4115 565 4167
rect 617 4115 623 4167
rect 726 4110 732 4162
rect 784 4110 790 4162
rect 1151 4109 1157 4161
rect 1209 4109 1215 4161
rect 1794 4122 1800 4174
rect 1852 4122 1858 4174
rect 3042 4122 3048 4174
rect 3100 4122 3106 4174
rect 559 3733 565 3785
rect 617 3733 623 3785
rect 726 3738 732 3790
rect 784 3738 790 3790
rect 1151 3739 1157 3791
rect 1209 3739 1215 3791
rect 1794 3726 1800 3778
rect 1852 3726 1858 3778
rect 3042 3726 3048 3778
rect 3100 3726 3106 3778
rect 559 3325 565 3377
rect 617 3325 623 3377
rect 726 3320 732 3372
rect 784 3320 790 3372
rect 1151 3319 1157 3371
rect 1209 3319 1215 3371
rect 1794 3332 1800 3384
rect 1852 3332 1858 3384
rect 3042 3332 3048 3384
rect 3100 3332 3106 3384
rect 559 2943 565 2995
rect 617 2943 623 2995
rect 726 2948 732 3000
rect 784 2948 790 3000
rect 1151 2949 1157 3001
rect 1209 2949 1215 3001
rect 1794 2936 1800 2988
rect 1852 2936 1858 2988
rect 3042 2936 3048 2988
rect 3100 2936 3106 2988
rect 559 2535 565 2587
rect 617 2535 623 2587
rect 726 2530 732 2582
rect 784 2530 790 2582
rect 1151 2529 1157 2581
rect 1209 2529 1215 2581
rect 1794 2542 1800 2594
rect 1852 2542 1858 2594
rect 3042 2542 3048 2594
rect 3100 2542 3106 2594
rect 559 2153 565 2205
rect 617 2153 623 2205
rect 726 2158 732 2210
rect 784 2158 790 2210
rect 1151 2159 1157 2211
rect 1209 2159 1215 2211
rect 1794 2146 1800 2198
rect 1852 2146 1858 2198
rect 3042 2146 3048 2198
rect 3100 2146 3106 2198
rect 559 1745 565 1797
rect 617 1745 623 1797
rect 726 1740 732 1792
rect 784 1740 790 1792
rect 1151 1739 1157 1791
rect 1209 1739 1215 1791
rect 1794 1752 1800 1804
rect 1852 1752 1858 1804
rect 3042 1752 3048 1804
rect 3100 1752 3106 1804
rect 559 1363 565 1415
rect 617 1363 623 1415
rect 726 1368 732 1420
rect 784 1368 790 1420
rect 1151 1369 1157 1421
rect 1209 1369 1215 1421
rect 1794 1356 1800 1408
rect 1852 1356 1858 1408
rect 3042 1356 3048 1408
rect 3100 1356 3106 1408
rect 559 955 565 1007
rect 617 955 623 1007
rect 726 950 732 1002
rect 784 950 790 1002
rect 1151 949 1157 1001
rect 1209 949 1215 1001
rect 1794 962 1800 1014
rect 1852 962 1858 1014
rect 3042 962 3048 1014
rect 3100 962 3106 1014
rect 559 573 565 625
rect 617 573 623 625
rect 726 578 732 630
rect 784 578 790 630
rect 1151 579 1157 631
rect 1209 579 1215 631
rect 1794 566 1800 618
rect 1852 566 1858 618
rect 3042 566 3048 618
rect 3100 566 3106 618
rect 559 165 565 217
rect 617 165 623 217
rect 726 160 732 212
rect 784 160 790 212
rect 1151 159 1157 211
rect 1209 159 1215 211
rect 1794 172 1800 224
rect 1852 172 1858 224
rect 3042 172 3048 224
rect 3100 172 3106 224
<< via1 >>
rect 565 25106 617 25115
rect 565 25072 574 25106
rect 574 25072 608 25106
rect 608 25072 617 25106
rect 565 25063 617 25072
rect 732 25068 784 25120
rect 1157 25069 1209 25121
rect 1800 25056 1852 25108
rect 3048 25056 3100 25108
rect 565 24698 617 24707
rect 565 24664 574 24698
rect 574 24664 608 24698
rect 608 24664 617 24698
rect 565 24655 617 24664
rect 732 24650 784 24702
rect 1157 24649 1209 24701
rect 1800 24662 1852 24714
rect 3048 24662 3100 24714
rect 565 24316 617 24325
rect 565 24282 574 24316
rect 574 24282 608 24316
rect 608 24282 617 24316
rect 565 24273 617 24282
rect 732 24278 784 24330
rect 1157 24279 1209 24331
rect 1800 24266 1852 24318
rect 3048 24266 3100 24318
rect 565 23908 617 23917
rect 565 23874 574 23908
rect 574 23874 608 23908
rect 608 23874 617 23908
rect 565 23865 617 23874
rect 732 23860 784 23912
rect 1157 23859 1209 23911
rect 1800 23872 1852 23924
rect 3048 23872 3100 23924
rect 565 23526 617 23535
rect 565 23492 574 23526
rect 574 23492 608 23526
rect 608 23492 617 23526
rect 565 23483 617 23492
rect 732 23488 784 23540
rect 1157 23489 1209 23541
rect 1800 23476 1852 23528
rect 3048 23476 3100 23528
rect 565 23118 617 23127
rect 565 23084 574 23118
rect 574 23084 608 23118
rect 608 23084 617 23118
rect 565 23075 617 23084
rect 732 23070 784 23122
rect 1157 23069 1209 23121
rect 1800 23082 1852 23134
rect 3048 23082 3100 23134
rect 565 22736 617 22745
rect 565 22702 574 22736
rect 574 22702 608 22736
rect 608 22702 617 22736
rect 565 22693 617 22702
rect 732 22698 784 22750
rect 1157 22699 1209 22751
rect 1800 22686 1852 22738
rect 3048 22686 3100 22738
rect 565 22328 617 22337
rect 565 22294 574 22328
rect 574 22294 608 22328
rect 608 22294 617 22328
rect 565 22285 617 22294
rect 732 22280 784 22332
rect 1157 22279 1209 22331
rect 1800 22292 1852 22344
rect 3048 22292 3100 22344
rect 565 21946 617 21955
rect 565 21912 574 21946
rect 574 21912 608 21946
rect 608 21912 617 21946
rect 565 21903 617 21912
rect 732 21908 784 21960
rect 1157 21909 1209 21961
rect 1800 21896 1852 21948
rect 3048 21896 3100 21948
rect 565 21538 617 21547
rect 565 21504 574 21538
rect 574 21504 608 21538
rect 608 21504 617 21538
rect 565 21495 617 21504
rect 732 21490 784 21542
rect 1157 21489 1209 21541
rect 1800 21502 1852 21554
rect 3048 21502 3100 21554
rect 565 21156 617 21165
rect 565 21122 574 21156
rect 574 21122 608 21156
rect 608 21122 617 21156
rect 565 21113 617 21122
rect 732 21118 784 21170
rect 1157 21119 1209 21171
rect 1800 21106 1852 21158
rect 3048 21106 3100 21158
rect 565 20748 617 20757
rect 565 20714 574 20748
rect 574 20714 608 20748
rect 608 20714 617 20748
rect 565 20705 617 20714
rect 732 20700 784 20752
rect 1157 20699 1209 20751
rect 1800 20712 1852 20764
rect 3048 20712 3100 20764
rect 565 20366 617 20375
rect 565 20332 574 20366
rect 574 20332 608 20366
rect 608 20332 617 20366
rect 565 20323 617 20332
rect 732 20328 784 20380
rect 1157 20329 1209 20381
rect 1800 20316 1852 20368
rect 3048 20316 3100 20368
rect 565 19958 617 19967
rect 565 19924 574 19958
rect 574 19924 608 19958
rect 608 19924 617 19958
rect 565 19915 617 19924
rect 732 19910 784 19962
rect 1157 19909 1209 19961
rect 1800 19922 1852 19974
rect 3048 19922 3100 19974
rect 565 19576 617 19585
rect 565 19542 574 19576
rect 574 19542 608 19576
rect 608 19542 617 19576
rect 565 19533 617 19542
rect 732 19538 784 19590
rect 1157 19539 1209 19591
rect 1800 19526 1852 19578
rect 3048 19526 3100 19578
rect 565 19168 617 19177
rect 565 19134 574 19168
rect 574 19134 608 19168
rect 608 19134 617 19168
rect 565 19125 617 19134
rect 732 19120 784 19172
rect 1157 19119 1209 19171
rect 1800 19132 1852 19184
rect 3048 19132 3100 19184
rect 565 18786 617 18795
rect 565 18752 574 18786
rect 574 18752 608 18786
rect 608 18752 617 18786
rect 565 18743 617 18752
rect 732 18748 784 18800
rect 1157 18749 1209 18801
rect 1800 18736 1852 18788
rect 3048 18736 3100 18788
rect 565 18378 617 18387
rect 565 18344 574 18378
rect 574 18344 608 18378
rect 608 18344 617 18378
rect 565 18335 617 18344
rect 732 18330 784 18382
rect 1157 18329 1209 18381
rect 1800 18342 1852 18394
rect 3048 18342 3100 18394
rect 565 17996 617 18005
rect 565 17962 574 17996
rect 574 17962 608 17996
rect 608 17962 617 17996
rect 565 17953 617 17962
rect 732 17958 784 18010
rect 1157 17959 1209 18011
rect 1800 17946 1852 17998
rect 3048 17946 3100 17998
rect 565 17588 617 17597
rect 565 17554 574 17588
rect 574 17554 608 17588
rect 608 17554 617 17588
rect 565 17545 617 17554
rect 732 17540 784 17592
rect 1157 17539 1209 17591
rect 1800 17552 1852 17604
rect 3048 17552 3100 17604
rect 565 17206 617 17215
rect 565 17172 574 17206
rect 574 17172 608 17206
rect 608 17172 617 17206
rect 565 17163 617 17172
rect 732 17168 784 17220
rect 1157 17169 1209 17221
rect 1800 17156 1852 17208
rect 3048 17156 3100 17208
rect 565 16798 617 16807
rect 565 16764 574 16798
rect 574 16764 608 16798
rect 608 16764 617 16798
rect 565 16755 617 16764
rect 732 16750 784 16802
rect 1157 16749 1209 16801
rect 1800 16762 1852 16814
rect 3048 16762 3100 16814
rect 565 16416 617 16425
rect 565 16382 574 16416
rect 574 16382 608 16416
rect 608 16382 617 16416
rect 565 16373 617 16382
rect 732 16378 784 16430
rect 1157 16379 1209 16431
rect 1800 16366 1852 16418
rect 3048 16366 3100 16418
rect 565 16008 617 16017
rect 565 15974 574 16008
rect 574 15974 608 16008
rect 608 15974 617 16008
rect 565 15965 617 15974
rect 732 15960 784 16012
rect 1157 15959 1209 16011
rect 1800 15972 1852 16024
rect 3048 15972 3100 16024
rect 565 15626 617 15635
rect 565 15592 574 15626
rect 574 15592 608 15626
rect 608 15592 617 15626
rect 565 15583 617 15592
rect 732 15588 784 15640
rect 1157 15589 1209 15641
rect 1800 15576 1852 15628
rect 3048 15576 3100 15628
rect 565 15218 617 15227
rect 565 15184 574 15218
rect 574 15184 608 15218
rect 608 15184 617 15218
rect 565 15175 617 15184
rect 732 15170 784 15222
rect 1157 15169 1209 15221
rect 1800 15182 1852 15234
rect 3048 15182 3100 15234
rect 565 14836 617 14845
rect 565 14802 574 14836
rect 574 14802 608 14836
rect 608 14802 617 14836
rect 565 14793 617 14802
rect 732 14798 784 14850
rect 1157 14799 1209 14851
rect 1800 14786 1852 14838
rect 3048 14786 3100 14838
rect 565 14428 617 14437
rect 565 14394 574 14428
rect 574 14394 608 14428
rect 608 14394 617 14428
rect 565 14385 617 14394
rect 732 14380 784 14432
rect 1157 14379 1209 14431
rect 1800 14392 1852 14444
rect 3048 14392 3100 14444
rect 565 14046 617 14055
rect 565 14012 574 14046
rect 574 14012 608 14046
rect 608 14012 617 14046
rect 565 14003 617 14012
rect 732 14008 784 14060
rect 1157 14009 1209 14061
rect 1800 13996 1852 14048
rect 3048 13996 3100 14048
rect 565 13638 617 13647
rect 565 13604 574 13638
rect 574 13604 608 13638
rect 608 13604 617 13638
rect 565 13595 617 13604
rect 732 13590 784 13642
rect 1157 13589 1209 13641
rect 1800 13602 1852 13654
rect 3048 13602 3100 13654
rect 565 13256 617 13265
rect 565 13222 574 13256
rect 574 13222 608 13256
rect 608 13222 617 13256
rect 565 13213 617 13222
rect 732 13218 784 13270
rect 1157 13219 1209 13271
rect 1800 13206 1852 13258
rect 3048 13206 3100 13258
rect 565 12848 617 12857
rect 565 12814 574 12848
rect 574 12814 608 12848
rect 608 12814 617 12848
rect 565 12805 617 12814
rect 732 12800 784 12852
rect 1157 12799 1209 12851
rect 1800 12812 1852 12864
rect 3048 12812 3100 12864
rect 565 12466 617 12475
rect 565 12432 574 12466
rect 574 12432 608 12466
rect 608 12432 617 12466
rect 565 12423 617 12432
rect 732 12428 784 12480
rect 1157 12429 1209 12481
rect 1800 12416 1852 12468
rect 3048 12416 3100 12468
rect 565 12058 617 12067
rect 565 12024 574 12058
rect 574 12024 608 12058
rect 608 12024 617 12058
rect 565 12015 617 12024
rect 732 12010 784 12062
rect 1157 12009 1209 12061
rect 1800 12022 1852 12074
rect 3048 12022 3100 12074
rect 565 11676 617 11685
rect 565 11642 574 11676
rect 574 11642 608 11676
rect 608 11642 617 11676
rect 565 11633 617 11642
rect 732 11638 784 11690
rect 1157 11639 1209 11691
rect 1800 11626 1852 11678
rect 3048 11626 3100 11678
rect 565 11268 617 11277
rect 565 11234 574 11268
rect 574 11234 608 11268
rect 608 11234 617 11268
rect 565 11225 617 11234
rect 732 11220 784 11272
rect 1157 11219 1209 11271
rect 1800 11232 1852 11284
rect 3048 11232 3100 11284
rect 565 10886 617 10895
rect 565 10852 574 10886
rect 574 10852 608 10886
rect 608 10852 617 10886
rect 565 10843 617 10852
rect 732 10848 784 10900
rect 1157 10849 1209 10901
rect 1800 10836 1852 10888
rect 3048 10836 3100 10888
rect 565 10478 617 10487
rect 565 10444 574 10478
rect 574 10444 608 10478
rect 608 10444 617 10478
rect 565 10435 617 10444
rect 732 10430 784 10482
rect 1157 10429 1209 10481
rect 1800 10442 1852 10494
rect 3048 10442 3100 10494
rect 565 10096 617 10105
rect 565 10062 574 10096
rect 574 10062 608 10096
rect 608 10062 617 10096
rect 565 10053 617 10062
rect 732 10058 784 10110
rect 1157 10059 1209 10111
rect 1800 10046 1852 10098
rect 3048 10046 3100 10098
rect 565 9688 617 9697
rect 565 9654 574 9688
rect 574 9654 608 9688
rect 608 9654 617 9688
rect 565 9645 617 9654
rect 732 9640 784 9692
rect 1157 9639 1209 9691
rect 1800 9652 1852 9704
rect 3048 9652 3100 9704
rect 565 9306 617 9315
rect 565 9272 574 9306
rect 574 9272 608 9306
rect 608 9272 617 9306
rect 565 9263 617 9272
rect 732 9268 784 9320
rect 1157 9269 1209 9321
rect 1800 9256 1852 9308
rect 3048 9256 3100 9308
rect 565 8898 617 8907
rect 565 8864 574 8898
rect 574 8864 608 8898
rect 608 8864 617 8898
rect 565 8855 617 8864
rect 732 8850 784 8902
rect 1157 8849 1209 8901
rect 1800 8862 1852 8914
rect 3048 8862 3100 8914
rect 565 8516 617 8525
rect 565 8482 574 8516
rect 574 8482 608 8516
rect 608 8482 617 8516
rect 565 8473 617 8482
rect 732 8478 784 8530
rect 1157 8479 1209 8531
rect 1800 8466 1852 8518
rect 3048 8466 3100 8518
rect 565 8108 617 8117
rect 565 8074 574 8108
rect 574 8074 608 8108
rect 608 8074 617 8108
rect 565 8065 617 8074
rect 732 8060 784 8112
rect 1157 8059 1209 8111
rect 1800 8072 1852 8124
rect 3048 8072 3100 8124
rect 565 7726 617 7735
rect 565 7692 574 7726
rect 574 7692 608 7726
rect 608 7692 617 7726
rect 565 7683 617 7692
rect 732 7688 784 7740
rect 1157 7689 1209 7741
rect 1800 7676 1852 7728
rect 3048 7676 3100 7728
rect 565 7318 617 7327
rect 565 7284 574 7318
rect 574 7284 608 7318
rect 608 7284 617 7318
rect 565 7275 617 7284
rect 732 7270 784 7322
rect 1157 7269 1209 7321
rect 1800 7282 1852 7334
rect 3048 7282 3100 7334
rect 565 6936 617 6945
rect 565 6902 574 6936
rect 574 6902 608 6936
rect 608 6902 617 6936
rect 565 6893 617 6902
rect 732 6898 784 6950
rect 1157 6899 1209 6951
rect 1800 6886 1852 6938
rect 3048 6886 3100 6938
rect 565 6528 617 6537
rect 565 6494 574 6528
rect 574 6494 608 6528
rect 608 6494 617 6528
rect 565 6485 617 6494
rect 732 6480 784 6532
rect 1157 6479 1209 6531
rect 1800 6492 1852 6544
rect 3048 6492 3100 6544
rect 565 6146 617 6155
rect 565 6112 574 6146
rect 574 6112 608 6146
rect 608 6112 617 6146
rect 565 6103 617 6112
rect 732 6108 784 6160
rect 1157 6109 1209 6161
rect 1800 6096 1852 6148
rect 3048 6096 3100 6148
rect 565 5738 617 5747
rect 565 5704 574 5738
rect 574 5704 608 5738
rect 608 5704 617 5738
rect 565 5695 617 5704
rect 732 5690 784 5742
rect 1157 5689 1209 5741
rect 1800 5702 1852 5754
rect 3048 5702 3100 5754
rect 565 5356 617 5365
rect 565 5322 574 5356
rect 574 5322 608 5356
rect 608 5322 617 5356
rect 565 5313 617 5322
rect 732 5318 784 5370
rect 1157 5319 1209 5371
rect 1800 5306 1852 5358
rect 3048 5306 3100 5358
rect 565 4948 617 4957
rect 565 4914 574 4948
rect 574 4914 608 4948
rect 608 4914 617 4948
rect 565 4905 617 4914
rect 732 4900 784 4952
rect 1157 4899 1209 4951
rect 1800 4912 1852 4964
rect 3048 4912 3100 4964
rect 565 4566 617 4575
rect 565 4532 574 4566
rect 574 4532 608 4566
rect 608 4532 617 4566
rect 565 4523 617 4532
rect 732 4528 784 4580
rect 1157 4529 1209 4581
rect 1800 4516 1852 4568
rect 3048 4516 3100 4568
rect 565 4158 617 4167
rect 565 4124 574 4158
rect 574 4124 608 4158
rect 608 4124 617 4158
rect 565 4115 617 4124
rect 732 4110 784 4162
rect 1157 4109 1209 4161
rect 1800 4122 1852 4174
rect 3048 4122 3100 4174
rect 565 3776 617 3785
rect 565 3742 574 3776
rect 574 3742 608 3776
rect 608 3742 617 3776
rect 565 3733 617 3742
rect 732 3738 784 3790
rect 1157 3739 1209 3791
rect 1800 3726 1852 3778
rect 3048 3726 3100 3778
rect 565 3368 617 3377
rect 565 3334 574 3368
rect 574 3334 608 3368
rect 608 3334 617 3368
rect 565 3325 617 3334
rect 732 3320 784 3372
rect 1157 3319 1209 3371
rect 1800 3332 1852 3384
rect 3048 3332 3100 3384
rect 565 2986 617 2995
rect 565 2952 574 2986
rect 574 2952 608 2986
rect 608 2952 617 2986
rect 565 2943 617 2952
rect 732 2948 784 3000
rect 1157 2949 1209 3001
rect 1800 2936 1852 2988
rect 3048 2936 3100 2988
rect 565 2578 617 2587
rect 565 2544 574 2578
rect 574 2544 608 2578
rect 608 2544 617 2578
rect 565 2535 617 2544
rect 732 2530 784 2582
rect 1157 2529 1209 2581
rect 1800 2542 1852 2594
rect 3048 2542 3100 2594
rect 565 2196 617 2205
rect 565 2162 574 2196
rect 574 2162 608 2196
rect 608 2162 617 2196
rect 565 2153 617 2162
rect 732 2158 784 2210
rect 1157 2159 1209 2211
rect 1800 2146 1852 2198
rect 3048 2146 3100 2198
rect 565 1788 617 1797
rect 565 1754 574 1788
rect 574 1754 608 1788
rect 608 1754 617 1788
rect 565 1745 617 1754
rect 732 1740 784 1792
rect 1157 1739 1209 1791
rect 1800 1752 1852 1804
rect 3048 1752 3100 1804
rect 565 1406 617 1415
rect 565 1372 574 1406
rect 574 1372 608 1406
rect 608 1372 617 1406
rect 565 1363 617 1372
rect 732 1368 784 1420
rect 1157 1369 1209 1421
rect 1800 1356 1852 1408
rect 3048 1356 3100 1408
rect 565 998 617 1007
rect 565 964 574 998
rect 574 964 608 998
rect 608 964 617 998
rect 565 955 617 964
rect 732 950 784 1002
rect 1157 949 1209 1001
rect 1800 962 1852 1014
rect 3048 962 3100 1014
rect 565 616 617 625
rect 565 582 574 616
rect 574 582 608 616
rect 608 582 617 616
rect 565 573 617 582
rect 732 578 784 630
rect 1157 579 1209 631
rect 1800 566 1852 618
rect 3048 566 3100 618
rect 565 208 617 217
rect 565 174 574 208
rect 574 174 608 208
rect 608 174 617 208
rect 565 165 617 174
rect 732 160 784 212
rect 1157 159 1209 211
rect 1800 172 1852 224
rect 3048 172 3100 224
<< metal2 >>
rect 577 25121 605 25280
rect 730 25122 786 25131
rect 565 25115 617 25121
rect 565 25057 617 25063
rect 730 25057 786 25066
rect 1155 25123 1211 25132
rect 1155 25058 1211 25067
rect 1798 25111 1854 25120
rect 577 24713 605 25057
rect 1798 25046 1854 25055
rect 3046 25111 3102 25120
rect 3046 25046 3102 25055
rect 1798 24715 1854 24724
rect 565 24707 617 24713
rect 565 24649 617 24655
rect 730 24704 786 24713
rect 577 24331 605 24649
rect 730 24639 786 24648
rect 1155 24703 1211 24712
rect 1798 24650 1854 24659
rect 3046 24715 3102 24724
rect 3046 24650 3102 24659
rect 1155 24638 1211 24647
rect 730 24332 786 24341
rect 565 24325 617 24331
rect 565 24267 617 24273
rect 730 24267 786 24276
rect 1155 24333 1211 24342
rect 1155 24268 1211 24277
rect 1798 24321 1854 24330
rect 577 23923 605 24267
rect 1798 24256 1854 24265
rect 3046 24321 3102 24330
rect 3046 24256 3102 24265
rect 1798 23925 1854 23934
rect 565 23917 617 23923
rect 565 23859 617 23865
rect 730 23914 786 23923
rect 577 23541 605 23859
rect 730 23849 786 23858
rect 1155 23913 1211 23922
rect 1798 23860 1854 23869
rect 3046 23925 3102 23934
rect 3046 23860 3102 23869
rect 1155 23848 1211 23857
rect 730 23542 786 23551
rect 565 23535 617 23541
rect 565 23477 617 23483
rect 730 23477 786 23486
rect 1155 23543 1211 23552
rect 1155 23478 1211 23487
rect 1798 23531 1854 23540
rect 577 23133 605 23477
rect 1798 23466 1854 23475
rect 3046 23531 3102 23540
rect 3046 23466 3102 23475
rect 1798 23135 1854 23144
rect 565 23127 617 23133
rect 565 23069 617 23075
rect 730 23124 786 23133
rect 577 22751 605 23069
rect 730 23059 786 23068
rect 1155 23123 1211 23132
rect 1798 23070 1854 23079
rect 3046 23135 3102 23144
rect 3046 23070 3102 23079
rect 1155 23058 1211 23067
rect 730 22752 786 22761
rect 565 22745 617 22751
rect 565 22687 617 22693
rect 730 22687 786 22696
rect 1155 22753 1211 22762
rect 1155 22688 1211 22697
rect 1798 22741 1854 22750
rect 577 22343 605 22687
rect 1798 22676 1854 22685
rect 3046 22741 3102 22750
rect 3046 22676 3102 22685
rect 1798 22345 1854 22354
rect 565 22337 617 22343
rect 565 22279 617 22285
rect 730 22334 786 22343
rect 577 21961 605 22279
rect 730 22269 786 22278
rect 1155 22333 1211 22342
rect 1798 22280 1854 22289
rect 3046 22345 3102 22354
rect 3046 22280 3102 22289
rect 1155 22268 1211 22277
rect 730 21962 786 21971
rect 565 21955 617 21961
rect 565 21897 617 21903
rect 730 21897 786 21906
rect 1155 21963 1211 21972
rect 1155 21898 1211 21907
rect 1798 21951 1854 21960
rect 577 21553 605 21897
rect 1798 21886 1854 21895
rect 3046 21951 3102 21960
rect 3046 21886 3102 21895
rect 1798 21555 1854 21564
rect 565 21547 617 21553
rect 565 21489 617 21495
rect 730 21544 786 21553
rect 577 21171 605 21489
rect 730 21479 786 21488
rect 1155 21543 1211 21552
rect 1798 21490 1854 21499
rect 3046 21555 3102 21564
rect 3046 21490 3102 21499
rect 1155 21478 1211 21487
rect 730 21172 786 21181
rect 565 21165 617 21171
rect 565 21107 617 21113
rect 730 21107 786 21116
rect 1155 21173 1211 21182
rect 1155 21108 1211 21117
rect 1798 21161 1854 21170
rect 577 20763 605 21107
rect 1798 21096 1854 21105
rect 3046 21161 3102 21170
rect 3046 21096 3102 21105
rect 1798 20765 1854 20774
rect 565 20757 617 20763
rect 565 20699 617 20705
rect 730 20754 786 20763
rect 577 20381 605 20699
rect 730 20689 786 20698
rect 1155 20753 1211 20762
rect 1798 20700 1854 20709
rect 3046 20765 3102 20774
rect 3046 20700 3102 20709
rect 1155 20688 1211 20697
rect 730 20382 786 20391
rect 565 20375 617 20381
rect 565 20317 617 20323
rect 730 20317 786 20326
rect 1155 20383 1211 20392
rect 1155 20318 1211 20327
rect 1798 20371 1854 20380
rect 577 19973 605 20317
rect 1798 20306 1854 20315
rect 3046 20371 3102 20380
rect 3046 20306 3102 20315
rect 1798 19975 1854 19984
rect 565 19967 617 19973
rect 565 19909 617 19915
rect 730 19964 786 19973
rect 577 19591 605 19909
rect 730 19899 786 19908
rect 1155 19963 1211 19972
rect 1798 19910 1854 19919
rect 3046 19975 3102 19984
rect 3046 19910 3102 19919
rect 1155 19898 1211 19907
rect 730 19592 786 19601
rect 565 19585 617 19591
rect 565 19527 617 19533
rect 730 19527 786 19536
rect 1155 19593 1211 19602
rect 1155 19528 1211 19537
rect 1798 19581 1854 19590
rect 577 19183 605 19527
rect 1798 19516 1854 19525
rect 3046 19581 3102 19590
rect 3046 19516 3102 19525
rect 1798 19185 1854 19194
rect 565 19177 617 19183
rect 565 19119 617 19125
rect 730 19174 786 19183
rect 577 18801 605 19119
rect 730 19109 786 19118
rect 1155 19173 1211 19182
rect 1798 19120 1854 19129
rect 3046 19185 3102 19194
rect 3046 19120 3102 19129
rect 1155 19108 1211 19117
rect 730 18802 786 18811
rect 565 18795 617 18801
rect 565 18737 617 18743
rect 730 18737 786 18746
rect 1155 18803 1211 18812
rect 1155 18738 1211 18747
rect 1798 18791 1854 18800
rect 577 18393 605 18737
rect 1798 18726 1854 18735
rect 3046 18791 3102 18800
rect 3046 18726 3102 18735
rect 1798 18395 1854 18404
rect 565 18387 617 18393
rect 565 18329 617 18335
rect 730 18384 786 18393
rect 577 18011 605 18329
rect 730 18319 786 18328
rect 1155 18383 1211 18392
rect 1798 18330 1854 18339
rect 3046 18395 3102 18404
rect 3046 18330 3102 18339
rect 1155 18318 1211 18327
rect 730 18012 786 18021
rect 565 18005 617 18011
rect 565 17947 617 17953
rect 730 17947 786 17956
rect 1155 18013 1211 18022
rect 1155 17948 1211 17957
rect 1798 18001 1854 18010
rect 577 17603 605 17947
rect 1798 17936 1854 17945
rect 3046 18001 3102 18010
rect 3046 17936 3102 17945
rect 1798 17605 1854 17614
rect 565 17597 617 17603
rect 565 17539 617 17545
rect 730 17594 786 17603
rect 577 17221 605 17539
rect 730 17529 786 17538
rect 1155 17593 1211 17602
rect 1798 17540 1854 17549
rect 3046 17605 3102 17614
rect 3046 17540 3102 17549
rect 1155 17528 1211 17537
rect 730 17222 786 17231
rect 565 17215 617 17221
rect 565 17157 617 17163
rect 730 17157 786 17166
rect 1155 17223 1211 17232
rect 1155 17158 1211 17167
rect 1798 17211 1854 17220
rect 577 16813 605 17157
rect 1798 17146 1854 17155
rect 3046 17211 3102 17220
rect 3046 17146 3102 17155
rect 1798 16815 1854 16824
rect 565 16807 617 16813
rect 565 16749 617 16755
rect 730 16804 786 16813
rect 577 16431 605 16749
rect 730 16739 786 16748
rect 1155 16803 1211 16812
rect 1798 16750 1854 16759
rect 3046 16815 3102 16824
rect 3046 16750 3102 16759
rect 1155 16738 1211 16747
rect 730 16432 786 16441
rect 565 16425 617 16431
rect 565 16367 617 16373
rect 730 16367 786 16376
rect 1155 16433 1211 16442
rect 1155 16368 1211 16377
rect 1798 16421 1854 16430
rect 577 16023 605 16367
rect 1798 16356 1854 16365
rect 3046 16421 3102 16430
rect 3046 16356 3102 16365
rect 1798 16025 1854 16034
rect 565 16017 617 16023
rect 565 15959 617 15965
rect 730 16014 786 16023
rect 577 15641 605 15959
rect 730 15949 786 15958
rect 1155 16013 1211 16022
rect 1798 15960 1854 15969
rect 3046 16025 3102 16034
rect 3046 15960 3102 15969
rect 1155 15948 1211 15957
rect 730 15642 786 15651
rect 565 15635 617 15641
rect 565 15577 617 15583
rect 730 15577 786 15586
rect 1155 15643 1211 15652
rect 1155 15578 1211 15587
rect 1798 15631 1854 15640
rect 577 15233 605 15577
rect 1798 15566 1854 15575
rect 3046 15631 3102 15640
rect 3046 15566 3102 15575
rect 1798 15235 1854 15244
rect 565 15227 617 15233
rect 565 15169 617 15175
rect 730 15224 786 15233
rect 577 14851 605 15169
rect 730 15159 786 15168
rect 1155 15223 1211 15232
rect 1798 15170 1854 15179
rect 3046 15235 3102 15244
rect 3046 15170 3102 15179
rect 1155 15158 1211 15167
rect 730 14852 786 14861
rect 565 14845 617 14851
rect 565 14787 617 14793
rect 730 14787 786 14796
rect 1155 14853 1211 14862
rect 1155 14788 1211 14797
rect 1798 14841 1854 14850
rect 577 14443 605 14787
rect 1798 14776 1854 14785
rect 3046 14841 3102 14850
rect 3046 14776 3102 14785
rect 1798 14445 1854 14454
rect 565 14437 617 14443
rect 565 14379 617 14385
rect 730 14434 786 14443
rect 577 14061 605 14379
rect 730 14369 786 14378
rect 1155 14433 1211 14442
rect 1798 14380 1854 14389
rect 3046 14445 3102 14454
rect 3046 14380 3102 14389
rect 1155 14368 1211 14377
rect 730 14062 786 14071
rect 565 14055 617 14061
rect 565 13997 617 14003
rect 730 13997 786 14006
rect 1155 14063 1211 14072
rect 1155 13998 1211 14007
rect 1798 14051 1854 14060
rect 577 13653 605 13997
rect 1798 13986 1854 13995
rect 3046 14051 3102 14060
rect 3046 13986 3102 13995
rect 1798 13655 1854 13664
rect 565 13647 617 13653
rect 565 13589 617 13595
rect 730 13644 786 13653
rect 577 13271 605 13589
rect 730 13579 786 13588
rect 1155 13643 1211 13652
rect 1798 13590 1854 13599
rect 3046 13655 3102 13664
rect 3046 13590 3102 13599
rect 1155 13578 1211 13587
rect 730 13272 786 13281
rect 565 13265 617 13271
rect 565 13207 617 13213
rect 730 13207 786 13216
rect 1155 13273 1211 13282
rect 1155 13208 1211 13217
rect 1798 13261 1854 13270
rect 577 12863 605 13207
rect 1798 13196 1854 13205
rect 3046 13261 3102 13270
rect 3046 13196 3102 13205
rect 1798 12865 1854 12874
rect 565 12857 617 12863
rect 565 12799 617 12805
rect 730 12854 786 12863
rect 577 12481 605 12799
rect 730 12789 786 12798
rect 1155 12853 1211 12862
rect 1798 12800 1854 12809
rect 3046 12865 3102 12874
rect 3046 12800 3102 12809
rect 1155 12788 1211 12797
rect 730 12482 786 12491
rect 565 12475 617 12481
rect 565 12417 617 12423
rect 730 12417 786 12426
rect 1155 12483 1211 12492
rect 1155 12418 1211 12427
rect 1798 12471 1854 12480
rect 577 12073 605 12417
rect 1798 12406 1854 12415
rect 3046 12471 3102 12480
rect 3046 12406 3102 12415
rect 1798 12075 1854 12084
rect 565 12067 617 12073
rect 565 12009 617 12015
rect 730 12064 786 12073
rect 577 11691 605 12009
rect 730 11999 786 12008
rect 1155 12063 1211 12072
rect 1798 12010 1854 12019
rect 3046 12075 3102 12084
rect 3046 12010 3102 12019
rect 1155 11998 1211 12007
rect 730 11692 786 11701
rect 565 11685 617 11691
rect 565 11627 617 11633
rect 730 11627 786 11636
rect 1155 11693 1211 11702
rect 1155 11628 1211 11637
rect 1798 11681 1854 11690
rect 577 11283 605 11627
rect 1798 11616 1854 11625
rect 3046 11681 3102 11690
rect 3046 11616 3102 11625
rect 1798 11285 1854 11294
rect 565 11277 617 11283
rect 565 11219 617 11225
rect 730 11274 786 11283
rect 577 10901 605 11219
rect 730 11209 786 11218
rect 1155 11273 1211 11282
rect 1798 11220 1854 11229
rect 3046 11285 3102 11294
rect 3046 11220 3102 11229
rect 1155 11208 1211 11217
rect 730 10902 786 10911
rect 565 10895 617 10901
rect 565 10837 617 10843
rect 730 10837 786 10846
rect 1155 10903 1211 10912
rect 1155 10838 1211 10847
rect 1798 10891 1854 10900
rect 577 10493 605 10837
rect 1798 10826 1854 10835
rect 3046 10891 3102 10900
rect 3046 10826 3102 10835
rect 1798 10495 1854 10504
rect 565 10487 617 10493
rect 565 10429 617 10435
rect 730 10484 786 10493
rect 577 10111 605 10429
rect 730 10419 786 10428
rect 1155 10483 1211 10492
rect 1798 10430 1854 10439
rect 3046 10495 3102 10504
rect 3046 10430 3102 10439
rect 1155 10418 1211 10427
rect 730 10112 786 10121
rect 565 10105 617 10111
rect 565 10047 617 10053
rect 730 10047 786 10056
rect 1155 10113 1211 10122
rect 1155 10048 1211 10057
rect 1798 10101 1854 10110
rect 577 9703 605 10047
rect 1798 10036 1854 10045
rect 3046 10101 3102 10110
rect 3046 10036 3102 10045
rect 1798 9705 1854 9714
rect 565 9697 617 9703
rect 565 9639 617 9645
rect 730 9694 786 9703
rect 577 9321 605 9639
rect 730 9629 786 9638
rect 1155 9693 1211 9702
rect 1798 9640 1854 9649
rect 3046 9705 3102 9714
rect 3046 9640 3102 9649
rect 1155 9628 1211 9637
rect 730 9322 786 9331
rect 565 9315 617 9321
rect 565 9257 617 9263
rect 730 9257 786 9266
rect 1155 9323 1211 9332
rect 1155 9258 1211 9267
rect 1798 9311 1854 9320
rect 577 8913 605 9257
rect 1798 9246 1854 9255
rect 3046 9311 3102 9320
rect 3046 9246 3102 9255
rect 1798 8915 1854 8924
rect 565 8907 617 8913
rect 565 8849 617 8855
rect 730 8904 786 8913
rect 577 8531 605 8849
rect 730 8839 786 8848
rect 1155 8903 1211 8912
rect 1798 8850 1854 8859
rect 3046 8915 3102 8924
rect 3046 8850 3102 8859
rect 1155 8838 1211 8847
rect 730 8532 786 8541
rect 565 8525 617 8531
rect 565 8467 617 8473
rect 730 8467 786 8476
rect 1155 8533 1211 8542
rect 1155 8468 1211 8477
rect 1798 8521 1854 8530
rect 577 8123 605 8467
rect 1798 8456 1854 8465
rect 3046 8521 3102 8530
rect 3046 8456 3102 8465
rect 1798 8125 1854 8134
rect 565 8117 617 8123
rect 565 8059 617 8065
rect 730 8114 786 8123
rect 577 7741 605 8059
rect 730 8049 786 8058
rect 1155 8113 1211 8122
rect 1798 8060 1854 8069
rect 3046 8125 3102 8134
rect 3046 8060 3102 8069
rect 1155 8048 1211 8057
rect 730 7742 786 7751
rect 565 7735 617 7741
rect 565 7677 617 7683
rect 730 7677 786 7686
rect 1155 7743 1211 7752
rect 1155 7678 1211 7687
rect 1798 7731 1854 7740
rect 577 7333 605 7677
rect 1798 7666 1854 7675
rect 3046 7731 3102 7740
rect 3046 7666 3102 7675
rect 1798 7335 1854 7344
rect 565 7327 617 7333
rect 565 7269 617 7275
rect 730 7324 786 7333
rect 577 6951 605 7269
rect 730 7259 786 7268
rect 1155 7323 1211 7332
rect 1798 7270 1854 7279
rect 3046 7335 3102 7344
rect 3046 7270 3102 7279
rect 1155 7258 1211 7267
rect 730 6952 786 6961
rect 565 6945 617 6951
rect 565 6887 617 6893
rect 730 6887 786 6896
rect 1155 6953 1211 6962
rect 1155 6888 1211 6897
rect 1798 6941 1854 6950
rect 577 6543 605 6887
rect 1798 6876 1854 6885
rect 3046 6941 3102 6950
rect 3046 6876 3102 6885
rect 1798 6545 1854 6554
rect 565 6537 617 6543
rect 565 6479 617 6485
rect 730 6534 786 6543
rect 577 6161 605 6479
rect 730 6469 786 6478
rect 1155 6533 1211 6542
rect 1798 6480 1854 6489
rect 3046 6545 3102 6554
rect 3046 6480 3102 6489
rect 1155 6468 1211 6477
rect 730 6162 786 6171
rect 565 6155 617 6161
rect 565 6097 617 6103
rect 730 6097 786 6106
rect 1155 6163 1211 6172
rect 1155 6098 1211 6107
rect 1798 6151 1854 6160
rect 577 5753 605 6097
rect 1798 6086 1854 6095
rect 3046 6151 3102 6160
rect 3046 6086 3102 6095
rect 1798 5755 1854 5764
rect 565 5747 617 5753
rect 565 5689 617 5695
rect 730 5744 786 5753
rect 577 5371 605 5689
rect 730 5679 786 5688
rect 1155 5743 1211 5752
rect 1798 5690 1854 5699
rect 3046 5755 3102 5764
rect 3046 5690 3102 5699
rect 1155 5678 1211 5687
rect 730 5372 786 5381
rect 565 5365 617 5371
rect 565 5307 617 5313
rect 730 5307 786 5316
rect 1155 5373 1211 5382
rect 1155 5308 1211 5317
rect 1798 5361 1854 5370
rect 577 4963 605 5307
rect 1798 5296 1854 5305
rect 3046 5361 3102 5370
rect 3046 5296 3102 5305
rect 1798 4965 1854 4974
rect 565 4957 617 4963
rect 565 4899 617 4905
rect 730 4954 786 4963
rect 577 4581 605 4899
rect 730 4889 786 4898
rect 1155 4953 1211 4962
rect 1798 4900 1854 4909
rect 3046 4965 3102 4974
rect 3046 4900 3102 4909
rect 1155 4888 1211 4897
rect 730 4582 786 4591
rect 565 4575 617 4581
rect 565 4517 617 4523
rect 730 4517 786 4526
rect 1155 4583 1211 4592
rect 1155 4518 1211 4527
rect 1798 4571 1854 4580
rect 577 4173 605 4517
rect 1798 4506 1854 4515
rect 3046 4571 3102 4580
rect 3046 4506 3102 4515
rect 1798 4175 1854 4184
rect 565 4167 617 4173
rect 565 4109 617 4115
rect 730 4164 786 4173
rect 577 3791 605 4109
rect 730 4099 786 4108
rect 1155 4163 1211 4172
rect 1798 4110 1854 4119
rect 3046 4175 3102 4184
rect 3046 4110 3102 4119
rect 1155 4098 1211 4107
rect 730 3792 786 3801
rect 565 3785 617 3791
rect 565 3727 617 3733
rect 730 3727 786 3736
rect 1155 3793 1211 3802
rect 1155 3728 1211 3737
rect 1798 3781 1854 3790
rect 577 3383 605 3727
rect 1798 3716 1854 3725
rect 3046 3781 3102 3790
rect 3046 3716 3102 3725
rect 1798 3385 1854 3394
rect 565 3377 617 3383
rect 565 3319 617 3325
rect 730 3374 786 3383
rect 577 3001 605 3319
rect 730 3309 786 3318
rect 1155 3373 1211 3382
rect 1798 3320 1854 3329
rect 3046 3385 3102 3394
rect 3046 3320 3102 3329
rect 1155 3308 1211 3317
rect 730 3002 786 3011
rect 565 2995 617 3001
rect 565 2937 617 2943
rect 730 2937 786 2946
rect 1155 3003 1211 3012
rect 1155 2938 1211 2947
rect 1798 2991 1854 3000
rect 577 2593 605 2937
rect 1798 2926 1854 2935
rect 3046 2991 3102 3000
rect 3046 2926 3102 2935
rect 1798 2595 1854 2604
rect 565 2587 617 2593
rect 565 2529 617 2535
rect 730 2584 786 2593
rect 577 2211 605 2529
rect 730 2519 786 2528
rect 1155 2583 1211 2592
rect 1798 2530 1854 2539
rect 3046 2595 3102 2604
rect 3046 2530 3102 2539
rect 1155 2518 1211 2527
rect 730 2212 786 2221
rect 565 2205 617 2211
rect 565 2147 617 2153
rect 730 2147 786 2156
rect 1155 2213 1211 2222
rect 1155 2148 1211 2157
rect 1798 2201 1854 2210
rect 577 1803 605 2147
rect 1798 2136 1854 2145
rect 3046 2201 3102 2210
rect 3046 2136 3102 2145
rect 1798 1805 1854 1814
rect 565 1797 617 1803
rect 565 1739 617 1745
rect 730 1794 786 1803
rect 577 1421 605 1739
rect 730 1729 786 1738
rect 1155 1793 1211 1802
rect 1798 1740 1854 1749
rect 3046 1805 3102 1814
rect 3046 1740 3102 1749
rect 1155 1728 1211 1737
rect 730 1422 786 1431
rect 565 1415 617 1421
rect 565 1357 617 1363
rect 730 1357 786 1366
rect 1155 1423 1211 1432
rect 1155 1358 1211 1367
rect 1798 1411 1854 1420
rect 577 1013 605 1357
rect 1798 1346 1854 1355
rect 3046 1411 3102 1420
rect 3046 1346 3102 1355
rect 1798 1015 1854 1024
rect 565 1007 617 1013
rect 565 949 617 955
rect 730 1004 786 1013
rect 577 631 605 949
rect 730 939 786 948
rect 1155 1003 1211 1012
rect 1798 950 1854 959
rect 3046 1015 3102 1024
rect 3046 950 3102 959
rect 1155 938 1211 947
rect 730 632 786 641
rect 565 625 617 631
rect 565 567 617 573
rect 730 567 786 576
rect 1155 633 1211 642
rect 1155 568 1211 577
rect 1798 621 1854 630
rect 577 223 605 567
rect 1798 556 1854 565
rect 3046 621 3102 630
rect 3046 556 3102 565
rect 1798 225 1854 234
rect 565 217 617 223
rect 565 159 617 165
rect 730 214 786 223
rect 577 0 605 159
rect 730 149 786 158
rect 1155 213 1211 222
rect 1798 160 1854 169
rect 3046 225 3102 234
rect 3046 160 3102 169
rect 1155 148 1211 157
<< via2 >>
rect 730 25120 786 25122
rect 730 25068 732 25120
rect 732 25068 784 25120
rect 784 25068 786 25120
rect 730 25066 786 25068
rect 1155 25121 1211 25123
rect 1155 25069 1157 25121
rect 1157 25069 1209 25121
rect 1209 25069 1211 25121
rect 1155 25067 1211 25069
rect 1798 25108 1854 25111
rect 1798 25056 1800 25108
rect 1800 25056 1852 25108
rect 1852 25056 1854 25108
rect 1798 25055 1854 25056
rect 3046 25108 3102 25111
rect 3046 25056 3048 25108
rect 3048 25056 3100 25108
rect 3100 25056 3102 25108
rect 3046 25055 3102 25056
rect 1798 24714 1854 24715
rect 730 24702 786 24704
rect 730 24650 732 24702
rect 732 24650 784 24702
rect 784 24650 786 24702
rect 730 24648 786 24650
rect 1155 24701 1211 24703
rect 1155 24649 1157 24701
rect 1157 24649 1209 24701
rect 1209 24649 1211 24701
rect 1798 24662 1800 24714
rect 1800 24662 1852 24714
rect 1852 24662 1854 24714
rect 1798 24659 1854 24662
rect 3046 24714 3102 24715
rect 3046 24662 3048 24714
rect 3048 24662 3100 24714
rect 3100 24662 3102 24714
rect 3046 24659 3102 24662
rect 1155 24647 1211 24649
rect 730 24330 786 24332
rect 730 24278 732 24330
rect 732 24278 784 24330
rect 784 24278 786 24330
rect 730 24276 786 24278
rect 1155 24331 1211 24333
rect 1155 24279 1157 24331
rect 1157 24279 1209 24331
rect 1209 24279 1211 24331
rect 1155 24277 1211 24279
rect 1798 24318 1854 24321
rect 1798 24266 1800 24318
rect 1800 24266 1852 24318
rect 1852 24266 1854 24318
rect 1798 24265 1854 24266
rect 3046 24318 3102 24321
rect 3046 24266 3048 24318
rect 3048 24266 3100 24318
rect 3100 24266 3102 24318
rect 3046 24265 3102 24266
rect 1798 23924 1854 23925
rect 730 23912 786 23914
rect 730 23860 732 23912
rect 732 23860 784 23912
rect 784 23860 786 23912
rect 730 23858 786 23860
rect 1155 23911 1211 23913
rect 1155 23859 1157 23911
rect 1157 23859 1209 23911
rect 1209 23859 1211 23911
rect 1798 23872 1800 23924
rect 1800 23872 1852 23924
rect 1852 23872 1854 23924
rect 1798 23869 1854 23872
rect 3046 23924 3102 23925
rect 3046 23872 3048 23924
rect 3048 23872 3100 23924
rect 3100 23872 3102 23924
rect 3046 23869 3102 23872
rect 1155 23857 1211 23859
rect 730 23540 786 23542
rect 730 23488 732 23540
rect 732 23488 784 23540
rect 784 23488 786 23540
rect 730 23486 786 23488
rect 1155 23541 1211 23543
rect 1155 23489 1157 23541
rect 1157 23489 1209 23541
rect 1209 23489 1211 23541
rect 1155 23487 1211 23489
rect 1798 23528 1854 23531
rect 1798 23476 1800 23528
rect 1800 23476 1852 23528
rect 1852 23476 1854 23528
rect 1798 23475 1854 23476
rect 3046 23528 3102 23531
rect 3046 23476 3048 23528
rect 3048 23476 3100 23528
rect 3100 23476 3102 23528
rect 3046 23475 3102 23476
rect 1798 23134 1854 23135
rect 730 23122 786 23124
rect 730 23070 732 23122
rect 732 23070 784 23122
rect 784 23070 786 23122
rect 730 23068 786 23070
rect 1155 23121 1211 23123
rect 1155 23069 1157 23121
rect 1157 23069 1209 23121
rect 1209 23069 1211 23121
rect 1798 23082 1800 23134
rect 1800 23082 1852 23134
rect 1852 23082 1854 23134
rect 1798 23079 1854 23082
rect 3046 23134 3102 23135
rect 3046 23082 3048 23134
rect 3048 23082 3100 23134
rect 3100 23082 3102 23134
rect 3046 23079 3102 23082
rect 1155 23067 1211 23069
rect 730 22750 786 22752
rect 730 22698 732 22750
rect 732 22698 784 22750
rect 784 22698 786 22750
rect 730 22696 786 22698
rect 1155 22751 1211 22753
rect 1155 22699 1157 22751
rect 1157 22699 1209 22751
rect 1209 22699 1211 22751
rect 1155 22697 1211 22699
rect 1798 22738 1854 22741
rect 1798 22686 1800 22738
rect 1800 22686 1852 22738
rect 1852 22686 1854 22738
rect 1798 22685 1854 22686
rect 3046 22738 3102 22741
rect 3046 22686 3048 22738
rect 3048 22686 3100 22738
rect 3100 22686 3102 22738
rect 3046 22685 3102 22686
rect 1798 22344 1854 22345
rect 730 22332 786 22334
rect 730 22280 732 22332
rect 732 22280 784 22332
rect 784 22280 786 22332
rect 730 22278 786 22280
rect 1155 22331 1211 22333
rect 1155 22279 1157 22331
rect 1157 22279 1209 22331
rect 1209 22279 1211 22331
rect 1798 22292 1800 22344
rect 1800 22292 1852 22344
rect 1852 22292 1854 22344
rect 1798 22289 1854 22292
rect 3046 22344 3102 22345
rect 3046 22292 3048 22344
rect 3048 22292 3100 22344
rect 3100 22292 3102 22344
rect 3046 22289 3102 22292
rect 1155 22277 1211 22279
rect 730 21960 786 21962
rect 730 21908 732 21960
rect 732 21908 784 21960
rect 784 21908 786 21960
rect 730 21906 786 21908
rect 1155 21961 1211 21963
rect 1155 21909 1157 21961
rect 1157 21909 1209 21961
rect 1209 21909 1211 21961
rect 1155 21907 1211 21909
rect 1798 21948 1854 21951
rect 1798 21896 1800 21948
rect 1800 21896 1852 21948
rect 1852 21896 1854 21948
rect 1798 21895 1854 21896
rect 3046 21948 3102 21951
rect 3046 21896 3048 21948
rect 3048 21896 3100 21948
rect 3100 21896 3102 21948
rect 3046 21895 3102 21896
rect 1798 21554 1854 21555
rect 730 21542 786 21544
rect 730 21490 732 21542
rect 732 21490 784 21542
rect 784 21490 786 21542
rect 730 21488 786 21490
rect 1155 21541 1211 21543
rect 1155 21489 1157 21541
rect 1157 21489 1209 21541
rect 1209 21489 1211 21541
rect 1798 21502 1800 21554
rect 1800 21502 1852 21554
rect 1852 21502 1854 21554
rect 1798 21499 1854 21502
rect 3046 21554 3102 21555
rect 3046 21502 3048 21554
rect 3048 21502 3100 21554
rect 3100 21502 3102 21554
rect 3046 21499 3102 21502
rect 1155 21487 1211 21489
rect 730 21170 786 21172
rect 730 21118 732 21170
rect 732 21118 784 21170
rect 784 21118 786 21170
rect 730 21116 786 21118
rect 1155 21171 1211 21173
rect 1155 21119 1157 21171
rect 1157 21119 1209 21171
rect 1209 21119 1211 21171
rect 1155 21117 1211 21119
rect 1798 21158 1854 21161
rect 1798 21106 1800 21158
rect 1800 21106 1852 21158
rect 1852 21106 1854 21158
rect 1798 21105 1854 21106
rect 3046 21158 3102 21161
rect 3046 21106 3048 21158
rect 3048 21106 3100 21158
rect 3100 21106 3102 21158
rect 3046 21105 3102 21106
rect 1798 20764 1854 20765
rect 730 20752 786 20754
rect 730 20700 732 20752
rect 732 20700 784 20752
rect 784 20700 786 20752
rect 730 20698 786 20700
rect 1155 20751 1211 20753
rect 1155 20699 1157 20751
rect 1157 20699 1209 20751
rect 1209 20699 1211 20751
rect 1798 20712 1800 20764
rect 1800 20712 1852 20764
rect 1852 20712 1854 20764
rect 1798 20709 1854 20712
rect 3046 20764 3102 20765
rect 3046 20712 3048 20764
rect 3048 20712 3100 20764
rect 3100 20712 3102 20764
rect 3046 20709 3102 20712
rect 1155 20697 1211 20699
rect 730 20380 786 20382
rect 730 20328 732 20380
rect 732 20328 784 20380
rect 784 20328 786 20380
rect 730 20326 786 20328
rect 1155 20381 1211 20383
rect 1155 20329 1157 20381
rect 1157 20329 1209 20381
rect 1209 20329 1211 20381
rect 1155 20327 1211 20329
rect 1798 20368 1854 20371
rect 1798 20316 1800 20368
rect 1800 20316 1852 20368
rect 1852 20316 1854 20368
rect 1798 20315 1854 20316
rect 3046 20368 3102 20371
rect 3046 20316 3048 20368
rect 3048 20316 3100 20368
rect 3100 20316 3102 20368
rect 3046 20315 3102 20316
rect 1798 19974 1854 19975
rect 730 19962 786 19964
rect 730 19910 732 19962
rect 732 19910 784 19962
rect 784 19910 786 19962
rect 730 19908 786 19910
rect 1155 19961 1211 19963
rect 1155 19909 1157 19961
rect 1157 19909 1209 19961
rect 1209 19909 1211 19961
rect 1798 19922 1800 19974
rect 1800 19922 1852 19974
rect 1852 19922 1854 19974
rect 1798 19919 1854 19922
rect 3046 19974 3102 19975
rect 3046 19922 3048 19974
rect 3048 19922 3100 19974
rect 3100 19922 3102 19974
rect 3046 19919 3102 19922
rect 1155 19907 1211 19909
rect 730 19590 786 19592
rect 730 19538 732 19590
rect 732 19538 784 19590
rect 784 19538 786 19590
rect 730 19536 786 19538
rect 1155 19591 1211 19593
rect 1155 19539 1157 19591
rect 1157 19539 1209 19591
rect 1209 19539 1211 19591
rect 1155 19537 1211 19539
rect 1798 19578 1854 19581
rect 1798 19526 1800 19578
rect 1800 19526 1852 19578
rect 1852 19526 1854 19578
rect 1798 19525 1854 19526
rect 3046 19578 3102 19581
rect 3046 19526 3048 19578
rect 3048 19526 3100 19578
rect 3100 19526 3102 19578
rect 3046 19525 3102 19526
rect 1798 19184 1854 19185
rect 730 19172 786 19174
rect 730 19120 732 19172
rect 732 19120 784 19172
rect 784 19120 786 19172
rect 730 19118 786 19120
rect 1155 19171 1211 19173
rect 1155 19119 1157 19171
rect 1157 19119 1209 19171
rect 1209 19119 1211 19171
rect 1798 19132 1800 19184
rect 1800 19132 1852 19184
rect 1852 19132 1854 19184
rect 1798 19129 1854 19132
rect 3046 19184 3102 19185
rect 3046 19132 3048 19184
rect 3048 19132 3100 19184
rect 3100 19132 3102 19184
rect 3046 19129 3102 19132
rect 1155 19117 1211 19119
rect 730 18800 786 18802
rect 730 18748 732 18800
rect 732 18748 784 18800
rect 784 18748 786 18800
rect 730 18746 786 18748
rect 1155 18801 1211 18803
rect 1155 18749 1157 18801
rect 1157 18749 1209 18801
rect 1209 18749 1211 18801
rect 1155 18747 1211 18749
rect 1798 18788 1854 18791
rect 1798 18736 1800 18788
rect 1800 18736 1852 18788
rect 1852 18736 1854 18788
rect 1798 18735 1854 18736
rect 3046 18788 3102 18791
rect 3046 18736 3048 18788
rect 3048 18736 3100 18788
rect 3100 18736 3102 18788
rect 3046 18735 3102 18736
rect 1798 18394 1854 18395
rect 730 18382 786 18384
rect 730 18330 732 18382
rect 732 18330 784 18382
rect 784 18330 786 18382
rect 730 18328 786 18330
rect 1155 18381 1211 18383
rect 1155 18329 1157 18381
rect 1157 18329 1209 18381
rect 1209 18329 1211 18381
rect 1798 18342 1800 18394
rect 1800 18342 1852 18394
rect 1852 18342 1854 18394
rect 1798 18339 1854 18342
rect 3046 18394 3102 18395
rect 3046 18342 3048 18394
rect 3048 18342 3100 18394
rect 3100 18342 3102 18394
rect 3046 18339 3102 18342
rect 1155 18327 1211 18329
rect 730 18010 786 18012
rect 730 17958 732 18010
rect 732 17958 784 18010
rect 784 17958 786 18010
rect 730 17956 786 17958
rect 1155 18011 1211 18013
rect 1155 17959 1157 18011
rect 1157 17959 1209 18011
rect 1209 17959 1211 18011
rect 1155 17957 1211 17959
rect 1798 17998 1854 18001
rect 1798 17946 1800 17998
rect 1800 17946 1852 17998
rect 1852 17946 1854 17998
rect 1798 17945 1854 17946
rect 3046 17998 3102 18001
rect 3046 17946 3048 17998
rect 3048 17946 3100 17998
rect 3100 17946 3102 17998
rect 3046 17945 3102 17946
rect 1798 17604 1854 17605
rect 730 17592 786 17594
rect 730 17540 732 17592
rect 732 17540 784 17592
rect 784 17540 786 17592
rect 730 17538 786 17540
rect 1155 17591 1211 17593
rect 1155 17539 1157 17591
rect 1157 17539 1209 17591
rect 1209 17539 1211 17591
rect 1798 17552 1800 17604
rect 1800 17552 1852 17604
rect 1852 17552 1854 17604
rect 1798 17549 1854 17552
rect 3046 17604 3102 17605
rect 3046 17552 3048 17604
rect 3048 17552 3100 17604
rect 3100 17552 3102 17604
rect 3046 17549 3102 17552
rect 1155 17537 1211 17539
rect 730 17220 786 17222
rect 730 17168 732 17220
rect 732 17168 784 17220
rect 784 17168 786 17220
rect 730 17166 786 17168
rect 1155 17221 1211 17223
rect 1155 17169 1157 17221
rect 1157 17169 1209 17221
rect 1209 17169 1211 17221
rect 1155 17167 1211 17169
rect 1798 17208 1854 17211
rect 1798 17156 1800 17208
rect 1800 17156 1852 17208
rect 1852 17156 1854 17208
rect 1798 17155 1854 17156
rect 3046 17208 3102 17211
rect 3046 17156 3048 17208
rect 3048 17156 3100 17208
rect 3100 17156 3102 17208
rect 3046 17155 3102 17156
rect 1798 16814 1854 16815
rect 730 16802 786 16804
rect 730 16750 732 16802
rect 732 16750 784 16802
rect 784 16750 786 16802
rect 730 16748 786 16750
rect 1155 16801 1211 16803
rect 1155 16749 1157 16801
rect 1157 16749 1209 16801
rect 1209 16749 1211 16801
rect 1798 16762 1800 16814
rect 1800 16762 1852 16814
rect 1852 16762 1854 16814
rect 1798 16759 1854 16762
rect 3046 16814 3102 16815
rect 3046 16762 3048 16814
rect 3048 16762 3100 16814
rect 3100 16762 3102 16814
rect 3046 16759 3102 16762
rect 1155 16747 1211 16749
rect 730 16430 786 16432
rect 730 16378 732 16430
rect 732 16378 784 16430
rect 784 16378 786 16430
rect 730 16376 786 16378
rect 1155 16431 1211 16433
rect 1155 16379 1157 16431
rect 1157 16379 1209 16431
rect 1209 16379 1211 16431
rect 1155 16377 1211 16379
rect 1798 16418 1854 16421
rect 1798 16366 1800 16418
rect 1800 16366 1852 16418
rect 1852 16366 1854 16418
rect 1798 16365 1854 16366
rect 3046 16418 3102 16421
rect 3046 16366 3048 16418
rect 3048 16366 3100 16418
rect 3100 16366 3102 16418
rect 3046 16365 3102 16366
rect 1798 16024 1854 16025
rect 730 16012 786 16014
rect 730 15960 732 16012
rect 732 15960 784 16012
rect 784 15960 786 16012
rect 730 15958 786 15960
rect 1155 16011 1211 16013
rect 1155 15959 1157 16011
rect 1157 15959 1209 16011
rect 1209 15959 1211 16011
rect 1798 15972 1800 16024
rect 1800 15972 1852 16024
rect 1852 15972 1854 16024
rect 1798 15969 1854 15972
rect 3046 16024 3102 16025
rect 3046 15972 3048 16024
rect 3048 15972 3100 16024
rect 3100 15972 3102 16024
rect 3046 15969 3102 15972
rect 1155 15957 1211 15959
rect 730 15640 786 15642
rect 730 15588 732 15640
rect 732 15588 784 15640
rect 784 15588 786 15640
rect 730 15586 786 15588
rect 1155 15641 1211 15643
rect 1155 15589 1157 15641
rect 1157 15589 1209 15641
rect 1209 15589 1211 15641
rect 1155 15587 1211 15589
rect 1798 15628 1854 15631
rect 1798 15576 1800 15628
rect 1800 15576 1852 15628
rect 1852 15576 1854 15628
rect 1798 15575 1854 15576
rect 3046 15628 3102 15631
rect 3046 15576 3048 15628
rect 3048 15576 3100 15628
rect 3100 15576 3102 15628
rect 3046 15575 3102 15576
rect 1798 15234 1854 15235
rect 730 15222 786 15224
rect 730 15170 732 15222
rect 732 15170 784 15222
rect 784 15170 786 15222
rect 730 15168 786 15170
rect 1155 15221 1211 15223
rect 1155 15169 1157 15221
rect 1157 15169 1209 15221
rect 1209 15169 1211 15221
rect 1798 15182 1800 15234
rect 1800 15182 1852 15234
rect 1852 15182 1854 15234
rect 1798 15179 1854 15182
rect 3046 15234 3102 15235
rect 3046 15182 3048 15234
rect 3048 15182 3100 15234
rect 3100 15182 3102 15234
rect 3046 15179 3102 15182
rect 1155 15167 1211 15169
rect 730 14850 786 14852
rect 730 14798 732 14850
rect 732 14798 784 14850
rect 784 14798 786 14850
rect 730 14796 786 14798
rect 1155 14851 1211 14853
rect 1155 14799 1157 14851
rect 1157 14799 1209 14851
rect 1209 14799 1211 14851
rect 1155 14797 1211 14799
rect 1798 14838 1854 14841
rect 1798 14786 1800 14838
rect 1800 14786 1852 14838
rect 1852 14786 1854 14838
rect 1798 14785 1854 14786
rect 3046 14838 3102 14841
rect 3046 14786 3048 14838
rect 3048 14786 3100 14838
rect 3100 14786 3102 14838
rect 3046 14785 3102 14786
rect 1798 14444 1854 14445
rect 730 14432 786 14434
rect 730 14380 732 14432
rect 732 14380 784 14432
rect 784 14380 786 14432
rect 730 14378 786 14380
rect 1155 14431 1211 14433
rect 1155 14379 1157 14431
rect 1157 14379 1209 14431
rect 1209 14379 1211 14431
rect 1798 14392 1800 14444
rect 1800 14392 1852 14444
rect 1852 14392 1854 14444
rect 1798 14389 1854 14392
rect 3046 14444 3102 14445
rect 3046 14392 3048 14444
rect 3048 14392 3100 14444
rect 3100 14392 3102 14444
rect 3046 14389 3102 14392
rect 1155 14377 1211 14379
rect 730 14060 786 14062
rect 730 14008 732 14060
rect 732 14008 784 14060
rect 784 14008 786 14060
rect 730 14006 786 14008
rect 1155 14061 1211 14063
rect 1155 14009 1157 14061
rect 1157 14009 1209 14061
rect 1209 14009 1211 14061
rect 1155 14007 1211 14009
rect 1798 14048 1854 14051
rect 1798 13996 1800 14048
rect 1800 13996 1852 14048
rect 1852 13996 1854 14048
rect 1798 13995 1854 13996
rect 3046 14048 3102 14051
rect 3046 13996 3048 14048
rect 3048 13996 3100 14048
rect 3100 13996 3102 14048
rect 3046 13995 3102 13996
rect 1798 13654 1854 13655
rect 730 13642 786 13644
rect 730 13590 732 13642
rect 732 13590 784 13642
rect 784 13590 786 13642
rect 730 13588 786 13590
rect 1155 13641 1211 13643
rect 1155 13589 1157 13641
rect 1157 13589 1209 13641
rect 1209 13589 1211 13641
rect 1798 13602 1800 13654
rect 1800 13602 1852 13654
rect 1852 13602 1854 13654
rect 1798 13599 1854 13602
rect 3046 13654 3102 13655
rect 3046 13602 3048 13654
rect 3048 13602 3100 13654
rect 3100 13602 3102 13654
rect 3046 13599 3102 13602
rect 1155 13587 1211 13589
rect 730 13270 786 13272
rect 730 13218 732 13270
rect 732 13218 784 13270
rect 784 13218 786 13270
rect 730 13216 786 13218
rect 1155 13271 1211 13273
rect 1155 13219 1157 13271
rect 1157 13219 1209 13271
rect 1209 13219 1211 13271
rect 1155 13217 1211 13219
rect 1798 13258 1854 13261
rect 1798 13206 1800 13258
rect 1800 13206 1852 13258
rect 1852 13206 1854 13258
rect 1798 13205 1854 13206
rect 3046 13258 3102 13261
rect 3046 13206 3048 13258
rect 3048 13206 3100 13258
rect 3100 13206 3102 13258
rect 3046 13205 3102 13206
rect 1798 12864 1854 12865
rect 730 12852 786 12854
rect 730 12800 732 12852
rect 732 12800 784 12852
rect 784 12800 786 12852
rect 730 12798 786 12800
rect 1155 12851 1211 12853
rect 1155 12799 1157 12851
rect 1157 12799 1209 12851
rect 1209 12799 1211 12851
rect 1798 12812 1800 12864
rect 1800 12812 1852 12864
rect 1852 12812 1854 12864
rect 1798 12809 1854 12812
rect 3046 12864 3102 12865
rect 3046 12812 3048 12864
rect 3048 12812 3100 12864
rect 3100 12812 3102 12864
rect 3046 12809 3102 12812
rect 1155 12797 1211 12799
rect 730 12480 786 12482
rect 730 12428 732 12480
rect 732 12428 784 12480
rect 784 12428 786 12480
rect 730 12426 786 12428
rect 1155 12481 1211 12483
rect 1155 12429 1157 12481
rect 1157 12429 1209 12481
rect 1209 12429 1211 12481
rect 1155 12427 1211 12429
rect 1798 12468 1854 12471
rect 1798 12416 1800 12468
rect 1800 12416 1852 12468
rect 1852 12416 1854 12468
rect 1798 12415 1854 12416
rect 3046 12468 3102 12471
rect 3046 12416 3048 12468
rect 3048 12416 3100 12468
rect 3100 12416 3102 12468
rect 3046 12415 3102 12416
rect 1798 12074 1854 12075
rect 730 12062 786 12064
rect 730 12010 732 12062
rect 732 12010 784 12062
rect 784 12010 786 12062
rect 730 12008 786 12010
rect 1155 12061 1211 12063
rect 1155 12009 1157 12061
rect 1157 12009 1209 12061
rect 1209 12009 1211 12061
rect 1798 12022 1800 12074
rect 1800 12022 1852 12074
rect 1852 12022 1854 12074
rect 1798 12019 1854 12022
rect 3046 12074 3102 12075
rect 3046 12022 3048 12074
rect 3048 12022 3100 12074
rect 3100 12022 3102 12074
rect 3046 12019 3102 12022
rect 1155 12007 1211 12009
rect 730 11690 786 11692
rect 730 11638 732 11690
rect 732 11638 784 11690
rect 784 11638 786 11690
rect 730 11636 786 11638
rect 1155 11691 1211 11693
rect 1155 11639 1157 11691
rect 1157 11639 1209 11691
rect 1209 11639 1211 11691
rect 1155 11637 1211 11639
rect 1798 11678 1854 11681
rect 1798 11626 1800 11678
rect 1800 11626 1852 11678
rect 1852 11626 1854 11678
rect 1798 11625 1854 11626
rect 3046 11678 3102 11681
rect 3046 11626 3048 11678
rect 3048 11626 3100 11678
rect 3100 11626 3102 11678
rect 3046 11625 3102 11626
rect 1798 11284 1854 11285
rect 730 11272 786 11274
rect 730 11220 732 11272
rect 732 11220 784 11272
rect 784 11220 786 11272
rect 730 11218 786 11220
rect 1155 11271 1211 11273
rect 1155 11219 1157 11271
rect 1157 11219 1209 11271
rect 1209 11219 1211 11271
rect 1798 11232 1800 11284
rect 1800 11232 1852 11284
rect 1852 11232 1854 11284
rect 1798 11229 1854 11232
rect 3046 11284 3102 11285
rect 3046 11232 3048 11284
rect 3048 11232 3100 11284
rect 3100 11232 3102 11284
rect 3046 11229 3102 11232
rect 1155 11217 1211 11219
rect 730 10900 786 10902
rect 730 10848 732 10900
rect 732 10848 784 10900
rect 784 10848 786 10900
rect 730 10846 786 10848
rect 1155 10901 1211 10903
rect 1155 10849 1157 10901
rect 1157 10849 1209 10901
rect 1209 10849 1211 10901
rect 1155 10847 1211 10849
rect 1798 10888 1854 10891
rect 1798 10836 1800 10888
rect 1800 10836 1852 10888
rect 1852 10836 1854 10888
rect 1798 10835 1854 10836
rect 3046 10888 3102 10891
rect 3046 10836 3048 10888
rect 3048 10836 3100 10888
rect 3100 10836 3102 10888
rect 3046 10835 3102 10836
rect 1798 10494 1854 10495
rect 730 10482 786 10484
rect 730 10430 732 10482
rect 732 10430 784 10482
rect 784 10430 786 10482
rect 730 10428 786 10430
rect 1155 10481 1211 10483
rect 1155 10429 1157 10481
rect 1157 10429 1209 10481
rect 1209 10429 1211 10481
rect 1798 10442 1800 10494
rect 1800 10442 1852 10494
rect 1852 10442 1854 10494
rect 1798 10439 1854 10442
rect 3046 10494 3102 10495
rect 3046 10442 3048 10494
rect 3048 10442 3100 10494
rect 3100 10442 3102 10494
rect 3046 10439 3102 10442
rect 1155 10427 1211 10429
rect 730 10110 786 10112
rect 730 10058 732 10110
rect 732 10058 784 10110
rect 784 10058 786 10110
rect 730 10056 786 10058
rect 1155 10111 1211 10113
rect 1155 10059 1157 10111
rect 1157 10059 1209 10111
rect 1209 10059 1211 10111
rect 1155 10057 1211 10059
rect 1798 10098 1854 10101
rect 1798 10046 1800 10098
rect 1800 10046 1852 10098
rect 1852 10046 1854 10098
rect 1798 10045 1854 10046
rect 3046 10098 3102 10101
rect 3046 10046 3048 10098
rect 3048 10046 3100 10098
rect 3100 10046 3102 10098
rect 3046 10045 3102 10046
rect 1798 9704 1854 9705
rect 730 9692 786 9694
rect 730 9640 732 9692
rect 732 9640 784 9692
rect 784 9640 786 9692
rect 730 9638 786 9640
rect 1155 9691 1211 9693
rect 1155 9639 1157 9691
rect 1157 9639 1209 9691
rect 1209 9639 1211 9691
rect 1798 9652 1800 9704
rect 1800 9652 1852 9704
rect 1852 9652 1854 9704
rect 1798 9649 1854 9652
rect 3046 9704 3102 9705
rect 3046 9652 3048 9704
rect 3048 9652 3100 9704
rect 3100 9652 3102 9704
rect 3046 9649 3102 9652
rect 1155 9637 1211 9639
rect 730 9320 786 9322
rect 730 9268 732 9320
rect 732 9268 784 9320
rect 784 9268 786 9320
rect 730 9266 786 9268
rect 1155 9321 1211 9323
rect 1155 9269 1157 9321
rect 1157 9269 1209 9321
rect 1209 9269 1211 9321
rect 1155 9267 1211 9269
rect 1798 9308 1854 9311
rect 1798 9256 1800 9308
rect 1800 9256 1852 9308
rect 1852 9256 1854 9308
rect 1798 9255 1854 9256
rect 3046 9308 3102 9311
rect 3046 9256 3048 9308
rect 3048 9256 3100 9308
rect 3100 9256 3102 9308
rect 3046 9255 3102 9256
rect 1798 8914 1854 8915
rect 730 8902 786 8904
rect 730 8850 732 8902
rect 732 8850 784 8902
rect 784 8850 786 8902
rect 730 8848 786 8850
rect 1155 8901 1211 8903
rect 1155 8849 1157 8901
rect 1157 8849 1209 8901
rect 1209 8849 1211 8901
rect 1798 8862 1800 8914
rect 1800 8862 1852 8914
rect 1852 8862 1854 8914
rect 1798 8859 1854 8862
rect 3046 8914 3102 8915
rect 3046 8862 3048 8914
rect 3048 8862 3100 8914
rect 3100 8862 3102 8914
rect 3046 8859 3102 8862
rect 1155 8847 1211 8849
rect 730 8530 786 8532
rect 730 8478 732 8530
rect 732 8478 784 8530
rect 784 8478 786 8530
rect 730 8476 786 8478
rect 1155 8531 1211 8533
rect 1155 8479 1157 8531
rect 1157 8479 1209 8531
rect 1209 8479 1211 8531
rect 1155 8477 1211 8479
rect 1798 8518 1854 8521
rect 1798 8466 1800 8518
rect 1800 8466 1852 8518
rect 1852 8466 1854 8518
rect 1798 8465 1854 8466
rect 3046 8518 3102 8521
rect 3046 8466 3048 8518
rect 3048 8466 3100 8518
rect 3100 8466 3102 8518
rect 3046 8465 3102 8466
rect 1798 8124 1854 8125
rect 730 8112 786 8114
rect 730 8060 732 8112
rect 732 8060 784 8112
rect 784 8060 786 8112
rect 730 8058 786 8060
rect 1155 8111 1211 8113
rect 1155 8059 1157 8111
rect 1157 8059 1209 8111
rect 1209 8059 1211 8111
rect 1798 8072 1800 8124
rect 1800 8072 1852 8124
rect 1852 8072 1854 8124
rect 1798 8069 1854 8072
rect 3046 8124 3102 8125
rect 3046 8072 3048 8124
rect 3048 8072 3100 8124
rect 3100 8072 3102 8124
rect 3046 8069 3102 8072
rect 1155 8057 1211 8059
rect 730 7740 786 7742
rect 730 7688 732 7740
rect 732 7688 784 7740
rect 784 7688 786 7740
rect 730 7686 786 7688
rect 1155 7741 1211 7743
rect 1155 7689 1157 7741
rect 1157 7689 1209 7741
rect 1209 7689 1211 7741
rect 1155 7687 1211 7689
rect 1798 7728 1854 7731
rect 1798 7676 1800 7728
rect 1800 7676 1852 7728
rect 1852 7676 1854 7728
rect 1798 7675 1854 7676
rect 3046 7728 3102 7731
rect 3046 7676 3048 7728
rect 3048 7676 3100 7728
rect 3100 7676 3102 7728
rect 3046 7675 3102 7676
rect 1798 7334 1854 7335
rect 730 7322 786 7324
rect 730 7270 732 7322
rect 732 7270 784 7322
rect 784 7270 786 7322
rect 730 7268 786 7270
rect 1155 7321 1211 7323
rect 1155 7269 1157 7321
rect 1157 7269 1209 7321
rect 1209 7269 1211 7321
rect 1798 7282 1800 7334
rect 1800 7282 1852 7334
rect 1852 7282 1854 7334
rect 1798 7279 1854 7282
rect 3046 7334 3102 7335
rect 3046 7282 3048 7334
rect 3048 7282 3100 7334
rect 3100 7282 3102 7334
rect 3046 7279 3102 7282
rect 1155 7267 1211 7269
rect 730 6950 786 6952
rect 730 6898 732 6950
rect 732 6898 784 6950
rect 784 6898 786 6950
rect 730 6896 786 6898
rect 1155 6951 1211 6953
rect 1155 6899 1157 6951
rect 1157 6899 1209 6951
rect 1209 6899 1211 6951
rect 1155 6897 1211 6899
rect 1798 6938 1854 6941
rect 1798 6886 1800 6938
rect 1800 6886 1852 6938
rect 1852 6886 1854 6938
rect 1798 6885 1854 6886
rect 3046 6938 3102 6941
rect 3046 6886 3048 6938
rect 3048 6886 3100 6938
rect 3100 6886 3102 6938
rect 3046 6885 3102 6886
rect 1798 6544 1854 6545
rect 730 6532 786 6534
rect 730 6480 732 6532
rect 732 6480 784 6532
rect 784 6480 786 6532
rect 730 6478 786 6480
rect 1155 6531 1211 6533
rect 1155 6479 1157 6531
rect 1157 6479 1209 6531
rect 1209 6479 1211 6531
rect 1798 6492 1800 6544
rect 1800 6492 1852 6544
rect 1852 6492 1854 6544
rect 1798 6489 1854 6492
rect 3046 6544 3102 6545
rect 3046 6492 3048 6544
rect 3048 6492 3100 6544
rect 3100 6492 3102 6544
rect 3046 6489 3102 6492
rect 1155 6477 1211 6479
rect 730 6160 786 6162
rect 730 6108 732 6160
rect 732 6108 784 6160
rect 784 6108 786 6160
rect 730 6106 786 6108
rect 1155 6161 1211 6163
rect 1155 6109 1157 6161
rect 1157 6109 1209 6161
rect 1209 6109 1211 6161
rect 1155 6107 1211 6109
rect 1798 6148 1854 6151
rect 1798 6096 1800 6148
rect 1800 6096 1852 6148
rect 1852 6096 1854 6148
rect 1798 6095 1854 6096
rect 3046 6148 3102 6151
rect 3046 6096 3048 6148
rect 3048 6096 3100 6148
rect 3100 6096 3102 6148
rect 3046 6095 3102 6096
rect 1798 5754 1854 5755
rect 730 5742 786 5744
rect 730 5690 732 5742
rect 732 5690 784 5742
rect 784 5690 786 5742
rect 730 5688 786 5690
rect 1155 5741 1211 5743
rect 1155 5689 1157 5741
rect 1157 5689 1209 5741
rect 1209 5689 1211 5741
rect 1798 5702 1800 5754
rect 1800 5702 1852 5754
rect 1852 5702 1854 5754
rect 1798 5699 1854 5702
rect 3046 5754 3102 5755
rect 3046 5702 3048 5754
rect 3048 5702 3100 5754
rect 3100 5702 3102 5754
rect 3046 5699 3102 5702
rect 1155 5687 1211 5689
rect 730 5370 786 5372
rect 730 5318 732 5370
rect 732 5318 784 5370
rect 784 5318 786 5370
rect 730 5316 786 5318
rect 1155 5371 1211 5373
rect 1155 5319 1157 5371
rect 1157 5319 1209 5371
rect 1209 5319 1211 5371
rect 1155 5317 1211 5319
rect 1798 5358 1854 5361
rect 1798 5306 1800 5358
rect 1800 5306 1852 5358
rect 1852 5306 1854 5358
rect 1798 5305 1854 5306
rect 3046 5358 3102 5361
rect 3046 5306 3048 5358
rect 3048 5306 3100 5358
rect 3100 5306 3102 5358
rect 3046 5305 3102 5306
rect 1798 4964 1854 4965
rect 730 4952 786 4954
rect 730 4900 732 4952
rect 732 4900 784 4952
rect 784 4900 786 4952
rect 730 4898 786 4900
rect 1155 4951 1211 4953
rect 1155 4899 1157 4951
rect 1157 4899 1209 4951
rect 1209 4899 1211 4951
rect 1798 4912 1800 4964
rect 1800 4912 1852 4964
rect 1852 4912 1854 4964
rect 1798 4909 1854 4912
rect 3046 4964 3102 4965
rect 3046 4912 3048 4964
rect 3048 4912 3100 4964
rect 3100 4912 3102 4964
rect 3046 4909 3102 4912
rect 1155 4897 1211 4899
rect 730 4580 786 4582
rect 730 4528 732 4580
rect 732 4528 784 4580
rect 784 4528 786 4580
rect 730 4526 786 4528
rect 1155 4581 1211 4583
rect 1155 4529 1157 4581
rect 1157 4529 1209 4581
rect 1209 4529 1211 4581
rect 1155 4527 1211 4529
rect 1798 4568 1854 4571
rect 1798 4516 1800 4568
rect 1800 4516 1852 4568
rect 1852 4516 1854 4568
rect 1798 4515 1854 4516
rect 3046 4568 3102 4571
rect 3046 4516 3048 4568
rect 3048 4516 3100 4568
rect 3100 4516 3102 4568
rect 3046 4515 3102 4516
rect 1798 4174 1854 4175
rect 730 4162 786 4164
rect 730 4110 732 4162
rect 732 4110 784 4162
rect 784 4110 786 4162
rect 730 4108 786 4110
rect 1155 4161 1211 4163
rect 1155 4109 1157 4161
rect 1157 4109 1209 4161
rect 1209 4109 1211 4161
rect 1798 4122 1800 4174
rect 1800 4122 1852 4174
rect 1852 4122 1854 4174
rect 1798 4119 1854 4122
rect 3046 4174 3102 4175
rect 3046 4122 3048 4174
rect 3048 4122 3100 4174
rect 3100 4122 3102 4174
rect 3046 4119 3102 4122
rect 1155 4107 1211 4109
rect 730 3790 786 3792
rect 730 3738 732 3790
rect 732 3738 784 3790
rect 784 3738 786 3790
rect 730 3736 786 3738
rect 1155 3791 1211 3793
rect 1155 3739 1157 3791
rect 1157 3739 1209 3791
rect 1209 3739 1211 3791
rect 1155 3737 1211 3739
rect 1798 3778 1854 3781
rect 1798 3726 1800 3778
rect 1800 3726 1852 3778
rect 1852 3726 1854 3778
rect 1798 3725 1854 3726
rect 3046 3778 3102 3781
rect 3046 3726 3048 3778
rect 3048 3726 3100 3778
rect 3100 3726 3102 3778
rect 3046 3725 3102 3726
rect 1798 3384 1854 3385
rect 730 3372 786 3374
rect 730 3320 732 3372
rect 732 3320 784 3372
rect 784 3320 786 3372
rect 730 3318 786 3320
rect 1155 3371 1211 3373
rect 1155 3319 1157 3371
rect 1157 3319 1209 3371
rect 1209 3319 1211 3371
rect 1798 3332 1800 3384
rect 1800 3332 1852 3384
rect 1852 3332 1854 3384
rect 1798 3329 1854 3332
rect 3046 3384 3102 3385
rect 3046 3332 3048 3384
rect 3048 3332 3100 3384
rect 3100 3332 3102 3384
rect 3046 3329 3102 3332
rect 1155 3317 1211 3319
rect 730 3000 786 3002
rect 730 2948 732 3000
rect 732 2948 784 3000
rect 784 2948 786 3000
rect 730 2946 786 2948
rect 1155 3001 1211 3003
rect 1155 2949 1157 3001
rect 1157 2949 1209 3001
rect 1209 2949 1211 3001
rect 1155 2947 1211 2949
rect 1798 2988 1854 2991
rect 1798 2936 1800 2988
rect 1800 2936 1852 2988
rect 1852 2936 1854 2988
rect 1798 2935 1854 2936
rect 3046 2988 3102 2991
rect 3046 2936 3048 2988
rect 3048 2936 3100 2988
rect 3100 2936 3102 2988
rect 3046 2935 3102 2936
rect 1798 2594 1854 2595
rect 730 2582 786 2584
rect 730 2530 732 2582
rect 732 2530 784 2582
rect 784 2530 786 2582
rect 730 2528 786 2530
rect 1155 2581 1211 2583
rect 1155 2529 1157 2581
rect 1157 2529 1209 2581
rect 1209 2529 1211 2581
rect 1798 2542 1800 2594
rect 1800 2542 1852 2594
rect 1852 2542 1854 2594
rect 1798 2539 1854 2542
rect 3046 2594 3102 2595
rect 3046 2542 3048 2594
rect 3048 2542 3100 2594
rect 3100 2542 3102 2594
rect 3046 2539 3102 2542
rect 1155 2527 1211 2529
rect 730 2210 786 2212
rect 730 2158 732 2210
rect 732 2158 784 2210
rect 784 2158 786 2210
rect 730 2156 786 2158
rect 1155 2211 1211 2213
rect 1155 2159 1157 2211
rect 1157 2159 1209 2211
rect 1209 2159 1211 2211
rect 1155 2157 1211 2159
rect 1798 2198 1854 2201
rect 1798 2146 1800 2198
rect 1800 2146 1852 2198
rect 1852 2146 1854 2198
rect 1798 2145 1854 2146
rect 3046 2198 3102 2201
rect 3046 2146 3048 2198
rect 3048 2146 3100 2198
rect 3100 2146 3102 2198
rect 3046 2145 3102 2146
rect 1798 1804 1854 1805
rect 730 1792 786 1794
rect 730 1740 732 1792
rect 732 1740 784 1792
rect 784 1740 786 1792
rect 730 1738 786 1740
rect 1155 1791 1211 1793
rect 1155 1739 1157 1791
rect 1157 1739 1209 1791
rect 1209 1739 1211 1791
rect 1798 1752 1800 1804
rect 1800 1752 1852 1804
rect 1852 1752 1854 1804
rect 1798 1749 1854 1752
rect 3046 1804 3102 1805
rect 3046 1752 3048 1804
rect 3048 1752 3100 1804
rect 3100 1752 3102 1804
rect 3046 1749 3102 1752
rect 1155 1737 1211 1739
rect 730 1420 786 1422
rect 730 1368 732 1420
rect 732 1368 784 1420
rect 784 1368 786 1420
rect 730 1366 786 1368
rect 1155 1421 1211 1423
rect 1155 1369 1157 1421
rect 1157 1369 1209 1421
rect 1209 1369 1211 1421
rect 1155 1367 1211 1369
rect 1798 1408 1854 1411
rect 1798 1356 1800 1408
rect 1800 1356 1852 1408
rect 1852 1356 1854 1408
rect 1798 1355 1854 1356
rect 3046 1408 3102 1411
rect 3046 1356 3048 1408
rect 3048 1356 3100 1408
rect 3100 1356 3102 1408
rect 3046 1355 3102 1356
rect 1798 1014 1854 1015
rect 730 1002 786 1004
rect 730 950 732 1002
rect 732 950 784 1002
rect 784 950 786 1002
rect 730 948 786 950
rect 1155 1001 1211 1003
rect 1155 949 1157 1001
rect 1157 949 1209 1001
rect 1209 949 1211 1001
rect 1798 962 1800 1014
rect 1800 962 1852 1014
rect 1852 962 1854 1014
rect 1798 959 1854 962
rect 3046 1014 3102 1015
rect 3046 962 3048 1014
rect 3048 962 3100 1014
rect 3100 962 3102 1014
rect 3046 959 3102 962
rect 1155 947 1211 949
rect 730 630 786 632
rect 730 578 732 630
rect 732 578 784 630
rect 784 578 786 630
rect 730 576 786 578
rect 1155 631 1211 633
rect 1155 579 1157 631
rect 1157 579 1209 631
rect 1209 579 1211 631
rect 1155 577 1211 579
rect 1798 618 1854 621
rect 1798 566 1800 618
rect 1800 566 1852 618
rect 1852 566 1854 618
rect 1798 565 1854 566
rect 3046 618 3102 621
rect 3046 566 3048 618
rect 3048 566 3100 618
rect 3100 566 3102 618
rect 3046 565 3102 566
rect 1798 224 1854 225
rect 730 212 786 214
rect 730 160 732 212
rect 732 160 784 212
rect 784 160 786 212
rect 730 158 786 160
rect 1155 211 1211 213
rect 1155 159 1157 211
rect 1157 159 1209 211
rect 1209 159 1211 211
rect 1798 172 1800 224
rect 1800 172 1852 224
rect 1852 172 1854 224
rect 1798 169 1854 172
rect 3046 224 3102 225
rect 3046 172 3048 224
rect 3048 172 3100 224
rect 3100 172 3102 224
rect 3046 169 3102 172
rect 1155 157 1211 159
<< metal3 >>
rect 1150 25127 1216 25128
rect 725 25126 791 25127
rect 683 25062 726 25126
rect 790 25062 833 25126
rect 1108 25063 1151 25127
rect 1215 25063 1258 25127
rect 1793 25115 1859 25116
rect 3041 25115 3107 25116
rect 1788 25114 1794 25115
rect 1150 25062 1216 25063
rect 725 25061 791 25062
rect 1751 25051 1794 25114
rect 1858 25114 1864 25115
rect 3036 25114 3042 25115
rect 1858 25051 1901 25114
rect 1751 25050 1901 25051
rect 2999 25051 3042 25114
rect 3106 25114 3112 25115
rect 3106 25051 3149 25114
rect 2999 25050 3149 25051
rect 1751 24719 1901 24720
rect 725 24708 791 24709
rect 683 24644 726 24708
rect 790 24644 833 24708
rect 1150 24707 1216 24708
rect 725 24643 791 24644
rect 1108 24643 1151 24707
rect 1215 24643 1258 24707
rect 1751 24656 1794 24719
rect 1788 24655 1794 24656
rect 1858 24656 1901 24719
rect 2999 24719 3149 24720
rect 2999 24656 3042 24719
rect 1858 24655 1864 24656
rect 3036 24655 3042 24656
rect 3106 24656 3149 24719
rect 3106 24655 3112 24656
rect 1793 24654 1859 24655
rect 3041 24654 3107 24655
rect 1150 24642 1216 24643
rect 1150 24337 1216 24338
rect 725 24336 791 24337
rect 683 24272 726 24336
rect 790 24272 833 24336
rect 1108 24273 1151 24337
rect 1215 24273 1258 24337
rect 1793 24325 1859 24326
rect 3041 24325 3107 24326
rect 1788 24324 1794 24325
rect 1150 24272 1216 24273
rect 725 24271 791 24272
rect 1751 24261 1794 24324
rect 1858 24324 1864 24325
rect 3036 24324 3042 24325
rect 1858 24261 1901 24324
rect 1751 24260 1901 24261
rect 2999 24261 3042 24324
rect 3106 24324 3112 24325
rect 3106 24261 3149 24324
rect 2999 24260 3149 24261
rect 1751 23929 1901 23930
rect 725 23918 791 23919
rect 683 23854 726 23918
rect 790 23854 833 23918
rect 1150 23917 1216 23918
rect 725 23853 791 23854
rect 1108 23853 1151 23917
rect 1215 23853 1258 23917
rect 1751 23866 1794 23929
rect 1788 23865 1794 23866
rect 1858 23866 1901 23929
rect 2999 23929 3149 23930
rect 2999 23866 3042 23929
rect 1858 23865 1864 23866
rect 3036 23865 3042 23866
rect 3106 23866 3149 23929
rect 3106 23865 3112 23866
rect 1793 23864 1859 23865
rect 3041 23864 3107 23865
rect 1150 23852 1216 23853
rect 1150 23547 1216 23548
rect 725 23546 791 23547
rect 683 23482 726 23546
rect 790 23482 833 23546
rect 1108 23483 1151 23547
rect 1215 23483 1258 23547
rect 1793 23535 1859 23536
rect 3041 23535 3107 23536
rect 1788 23534 1794 23535
rect 1150 23482 1216 23483
rect 725 23481 791 23482
rect 1751 23471 1794 23534
rect 1858 23534 1864 23535
rect 3036 23534 3042 23535
rect 1858 23471 1901 23534
rect 1751 23470 1901 23471
rect 2999 23471 3042 23534
rect 3106 23534 3112 23535
rect 3106 23471 3149 23534
rect 2999 23470 3149 23471
rect 1751 23139 1901 23140
rect 725 23128 791 23129
rect 683 23064 726 23128
rect 790 23064 833 23128
rect 1150 23127 1216 23128
rect 725 23063 791 23064
rect 1108 23063 1151 23127
rect 1215 23063 1258 23127
rect 1751 23076 1794 23139
rect 1788 23075 1794 23076
rect 1858 23076 1901 23139
rect 2999 23139 3149 23140
rect 2999 23076 3042 23139
rect 1858 23075 1864 23076
rect 3036 23075 3042 23076
rect 3106 23076 3149 23139
rect 3106 23075 3112 23076
rect 1793 23074 1859 23075
rect 3041 23074 3107 23075
rect 1150 23062 1216 23063
rect 1150 22757 1216 22758
rect 725 22756 791 22757
rect 683 22692 726 22756
rect 790 22692 833 22756
rect 1108 22693 1151 22757
rect 1215 22693 1258 22757
rect 1793 22745 1859 22746
rect 3041 22745 3107 22746
rect 1788 22744 1794 22745
rect 1150 22692 1216 22693
rect 725 22691 791 22692
rect 1751 22681 1794 22744
rect 1858 22744 1864 22745
rect 3036 22744 3042 22745
rect 1858 22681 1901 22744
rect 1751 22680 1901 22681
rect 2999 22681 3042 22744
rect 3106 22744 3112 22745
rect 3106 22681 3149 22744
rect 2999 22680 3149 22681
rect 1751 22349 1901 22350
rect 725 22338 791 22339
rect 683 22274 726 22338
rect 790 22274 833 22338
rect 1150 22337 1216 22338
rect 725 22273 791 22274
rect 1108 22273 1151 22337
rect 1215 22273 1258 22337
rect 1751 22286 1794 22349
rect 1788 22285 1794 22286
rect 1858 22286 1901 22349
rect 2999 22349 3149 22350
rect 2999 22286 3042 22349
rect 1858 22285 1864 22286
rect 3036 22285 3042 22286
rect 3106 22286 3149 22349
rect 3106 22285 3112 22286
rect 1793 22284 1859 22285
rect 3041 22284 3107 22285
rect 1150 22272 1216 22273
rect 1150 21967 1216 21968
rect 725 21966 791 21967
rect 683 21902 726 21966
rect 790 21902 833 21966
rect 1108 21903 1151 21967
rect 1215 21903 1258 21967
rect 1793 21955 1859 21956
rect 3041 21955 3107 21956
rect 1788 21954 1794 21955
rect 1150 21902 1216 21903
rect 725 21901 791 21902
rect 1751 21891 1794 21954
rect 1858 21954 1864 21955
rect 3036 21954 3042 21955
rect 1858 21891 1901 21954
rect 1751 21890 1901 21891
rect 2999 21891 3042 21954
rect 3106 21954 3112 21955
rect 3106 21891 3149 21954
rect 2999 21890 3149 21891
rect 1751 21559 1901 21560
rect 725 21548 791 21549
rect 683 21484 726 21548
rect 790 21484 833 21548
rect 1150 21547 1216 21548
rect 725 21483 791 21484
rect 1108 21483 1151 21547
rect 1215 21483 1258 21547
rect 1751 21496 1794 21559
rect 1788 21495 1794 21496
rect 1858 21496 1901 21559
rect 2999 21559 3149 21560
rect 2999 21496 3042 21559
rect 1858 21495 1864 21496
rect 3036 21495 3042 21496
rect 3106 21496 3149 21559
rect 3106 21495 3112 21496
rect 1793 21494 1859 21495
rect 3041 21494 3107 21495
rect 1150 21482 1216 21483
rect 1150 21177 1216 21178
rect 725 21176 791 21177
rect 683 21112 726 21176
rect 790 21112 833 21176
rect 1108 21113 1151 21177
rect 1215 21113 1258 21177
rect 1793 21165 1859 21166
rect 3041 21165 3107 21166
rect 1788 21164 1794 21165
rect 1150 21112 1216 21113
rect 725 21111 791 21112
rect 1751 21101 1794 21164
rect 1858 21164 1864 21165
rect 3036 21164 3042 21165
rect 1858 21101 1901 21164
rect 1751 21100 1901 21101
rect 2999 21101 3042 21164
rect 3106 21164 3112 21165
rect 3106 21101 3149 21164
rect 2999 21100 3149 21101
rect 1751 20769 1901 20770
rect 725 20758 791 20759
rect 683 20694 726 20758
rect 790 20694 833 20758
rect 1150 20757 1216 20758
rect 725 20693 791 20694
rect 1108 20693 1151 20757
rect 1215 20693 1258 20757
rect 1751 20706 1794 20769
rect 1788 20705 1794 20706
rect 1858 20706 1901 20769
rect 2999 20769 3149 20770
rect 2999 20706 3042 20769
rect 1858 20705 1864 20706
rect 3036 20705 3042 20706
rect 3106 20706 3149 20769
rect 3106 20705 3112 20706
rect 1793 20704 1859 20705
rect 3041 20704 3107 20705
rect 1150 20692 1216 20693
rect 1150 20387 1216 20388
rect 725 20386 791 20387
rect 683 20322 726 20386
rect 790 20322 833 20386
rect 1108 20323 1151 20387
rect 1215 20323 1258 20387
rect 1793 20375 1859 20376
rect 3041 20375 3107 20376
rect 1788 20374 1794 20375
rect 1150 20322 1216 20323
rect 725 20321 791 20322
rect 1751 20311 1794 20374
rect 1858 20374 1864 20375
rect 3036 20374 3042 20375
rect 1858 20311 1901 20374
rect 1751 20310 1901 20311
rect 2999 20311 3042 20374
rect 3106 20374 3112 20375
rect 3106 20311 3149 20374
rect 2999 20310 3149 20311
rect 1751 19979 1901 19980
rect 725 19968 791 19969
rect 683 19904 726 19968
rect 790 19904 833 19968
rect 1150 19967 1216 19968
rect 725 19903 791 19904
rect 1108 19903 1151 19967
rect 1215 19903 1258 19967
rect 1751 19916 1794 19979
rect 1788 19915 1794 19916
rect 1858 19916 1901 19979
rect 2999 19979 3149 19980
rect 2999 19916 3042 19979
rect 1858 19915 1864 19916
rect 3036 19915 3042 19916
rect 3106 19916 3149 19979
rect 3106 19915 3112 19916
rect 1793 19914 1859 19915
rect 3041 19914 3107 19915
rect 1150 19902 1216 19903
rect 1150 19597 1216 19598
rect 725 19596 791 19597
rect 683 19532 726 19596
rect 790 19532 833 19596
rect 1108 19533 1151 19597
rect 1215 19533 1258 19597
rect 1793 19585 1859 19586
rect 3041 19585 3107 19586
rect 1788 19584 1794 19585
rect 1150 19532 1216 19533
rect 725 19531 791 19532
rect 1751 19521 1794 19584
rect 1858 19584 1864 19585
rect 3036 19584 3042 19585
rect 1858 19521 1901 19584
rect 1751 19520 1901 19521
rect 2999 19521 3042 19584
rect 3106 19584 3112 19585
rect 3106 19521 3149 19584
rect 2999 19520 3149 19521
rect 1751 19189 1901 19190
rect 725 19178 791 19179
rect 683 19114 726 19178
rect 790 19114 833 19178
rect 1150 19177 1216 19178
rect 725 19113 791 19114
rect 1108 19113 1151 19177
rect 1215 19113 1258 19177
rect 1751 19126 1794 19189
rect 1788 19125 1794 19126
rect 1858 19126 1901 19189
rect 2999 19189 3149 19190
rect 2999 19126 3042 19189
rect 1858 19125 1864 19126
rect 3036 19125 3042 19126
rect 3106 19126 3149 19189
rect 3106 19125 3112 19126
rect 1793 19124 1859 19125
rect 3041 19124 3107 19125
rect 1150 19112 1216 19113
rect 1150 18807 1216 18808
rect 725 18806 791 18807
rect 683 18742 726 18806
rect 790 18742 833 18806
rect 1108 18743 1151 18807
rect 1215 18743 1258 18807
rect 1793 18795 1859 18796
rect 3041 18795 3107 18796
rect 1788 18794 1794 18795
rect 1150 18742 1216 18743
rect 725 18741 791 18742
rect 1751 18731 1794 18794
rect 1858 18794 1864 18795
rect 3036 18794 3042 18795
rect 1858 18731 1901 18794
rect 1751 18730 1901 18731
rect 2999 18731 3042 18794
rect 3106 18794 3112 18795
rect 3106 18731 3149 18794
rect 2999 18730 3149 18731
rect 1751 18399 1901 18400
rect 725 18388 791 18389
rect 683 18324 726 18388
rect 790 18324 833 18388
rect 1150 18387 1216 18388
rect 725 18323 791 18324
rect 1108 18323 1151 18387
rect 1215 18323 1258 18387
rect 1751 18336 1794 18399
rect 1788 18335 1794 18336
rect 1858 18336 1901 18399
rect 2999 18399 3149 18400
rect 2999 18336 3042 18399
rect 1858 18335 1864 18336
rect 3036 18335 3042 18336
rect 3106 18336 3149 18399
rect 3106 18335 3112 18336
rect 1793 18334 1859 18335
rect 3041 18334 3107 18335
rect 1150 18322 1216 18323
rect 1150 18017 1216 18018
rect 725 18016 791 18017
rect 683 17952 726 18016
rect 790 17952 833 18016
rect 1108 17953 1151 18017
rect 1215 17953 1258 18017
rect 1793 18005 1859 18006
rect 3041 18005 3107 18006
rect 1788 18004 1794 18005
rect 1150 17952 1216 17953
rect 725 17951 791 17952
rect 1751 17941 1794 18004
rect 1858 18004 1864 18005
rect 3036 18004 3042 18005
rect 1858 17941 1901 18004
rect 1751 17940 1901 17941
rect 2999 17941 3042 18004
rect 3106 18004 3112 18005
rect 3106 17941 3149 18004
rect 2999 17940 3149 17941
rect 1751 17609 1901 17610
rect 725 17598 791 17599
rect 683 17534 726 17598
rect 790 17534 833 17598
rect 1150 17597 1216 17598
rect 725 17533 791 17534
rect 1108 17533 1151 17597
rect 1215 17533 1258 17597
rect 1751 17546 1794 17609
rect 1788 17545 1794 17546
rect 1858 17546 1901 17609
rect 2999 17609 3149 17610
rect 2999 17546 3042 17609
rect 1858 17545 1864 17546
rect 3036 17545 3042 17546
rect 3106 17546 3149 17609
rect 3106 17545 3112 17546
rect 1793 17544 1859 17545
rect 3041 17544 3107 17545
rect 1150 17532 1216 17533
rect 1150 17227 1216 17228
rect 725 17226 791 17227
rect 683 17162 726 17226
rect 790 17162 833 17226
rect 1108 17163 1151 17227
rect 1215 17163 1258 17227
rect 1793 17215 1859 17216
rect 3041 17215 3107 17216
rect 1788 17214 1794 17215
rect 1150 17162 1216 17163
rect 725 17161 791 17162
rect 1751 17151 1794 17214
rect 1858 17214 1864 17215
rect 3036 17214 3042 17215
rect 1858 17151 1901 17214
rect 1751 17150 1901 17151
rect 2999 17151 3042 17214
rect 3106 17214 3112 17215
rect 3106 17151 3149 17214
rect 2999 17150 3149 17151
rect 1751 16819 1901 16820
rect 725 16808 791 16809
rect 683 16744 726 16808
rect 790 16744 833 16808
rect 1150 16807 1216 16808
rect 725 16743 791 16744
rect 1108 16743 1151 16807
rect 1215 16743 1258 16807
rect 1751 16756 1794 16819
rect 1788 16755 1794 16756
rect 1858 16756 1901 16819
rect 2999 16819 3149 16820
rect 2999 16756 3042 16819
rect 1858 16755 1864 16756
rect 3036 16755 3042 16756
rect 3106 16756 3149 16819
rect 3106 16755 3112 16756
rect 1793 16754 1859 16755
rect 3041 16754 3107 16755
rect 1150 16742 1216 16743
rect 1150 16437 1216 16438
rect 725 16436 791 16437
rect 683 16372 726 16436
rect 790 16372 833 16436
rect 1108 16373 1151 16437
rect 1215 16373 1258 16437
rect 1793 16425 1859 16426
rect 3041 16425 3107 16426
rect 1788 16424 1794 16425
rect 1150 16372 1216 16373
rect 725 16371 791 16372
rect 1751 16361 1794 16424
rect 1858 16424 1864 16425
rect 3036 16424 3042 16425
rect 1858 16361 1901 16424
rect 1751 16360 1901 16361
rect 2999 16361 3042 16424
rect 3106 16424 3112 16425
rect 3106 16361 3149 16424
rect 2999 16360 3149 16361
rect 1751 16029 1901 16030
rect 725 16018 791 16019
rect 683 15954 726 16018
rect 790 15954 833 16018
rect 1150 16017 1216 16018
rect 725 15953 791 15954
rect 1108 15953 1151 16017
rect 1215 15953 1258 16017
rect 1751 15966 1794 16029
rect 1788 15965 1794 15966
rect 1858 15966 1901 16029
rect 2999 16029 3149 16030
rect 2999 15966 3042 16029
rect 1858 15965 1864 15966
rect 3036 15965 3042 15966
rect 3106 15966 3149 16029
rect 3106 15965 3112 15966
rect 1793 15964 1859 15965
rect 3041 15964 3107 15965
rect 1150 15952 1216 15953
rect 1150 15647 1216 15648
rect 725 15646 791 15647
rect 683 15582 726 15646
rect 790 15582 833 15646
rect 1108 15583 1151 15647
rect 1215 15583 1258 15647
rect 1793 15635 1859 15636
rect 3041 15635 3107 15636
rect 1788 15634 1794 15635
rect 1150 15582 1216 15583
rect 725 15581 791 15582
rect 1751 15571 1794 15634
rect 1858 15634 1864 15635
rect 3036 15634 3042 15635
rect 1858 15571 1901 15634
rect 1751 15570 1901 15571
rect 2999 15571 3042 15634
rect 3106 15634 3112 15635
rect 3106 15571 3149 15634
rect 2999 15570 3149 15571
rect 1751 15239 1901 15240
rect 725 15228 791 15229
rect 683 15164 726 15228
rect 790 15164 833 15228
rect 1150 15227 1216 15228
rect 725 15163 791 15164
rect 1108 15163 1151 15227
rect 1215 15163 1258 15227
rect 1751 15176 1794 15239
rect 1788 15175 1794 15176
rect 1858 15176 1901 15239
rect 2999 15239 3149 15240
rect 2999 15176 3042 15239
rect 1858 15175 1864 15176
rect 3036 15175 3042 15176
rect 3106 15176 3149 15239
rect 3106 15175 3112 15176
rect 1793 15174 1859 15175
rect 3041 15174 3107 15175
rect 1150 15162 1216 15163
rect 1150 14857 1216 14858
rect 725 14856 791 14857
rect 683 14792 726 14856
rect 790 14792 833 14856
rect 1108 14793 1151 14857
rect 1215 14793 1258 14857
rect 1793 14845 1859 14846
rect 3041 14845 3107 14846
rect 1788 14844 1794 14845
rect 1150 14792 1216 14793
rect 725 14791 791 14792
rect 1751 14781 1794 14844
rect 1858 14844 1864 14845
rect 3036 14844 3042 14845
rect 1858 14781 1901 14844
rect 1751 14780 1901 14781
rect 2999 14781 3042 14844
rect 3106 14844 3112 14845
rect 3106 14781 3149 14844
rect 2999 14780 3149 14781
rect 1751 14449 1901 14450
rect 725 14438 791 14439
rect 683 14374 726 14438
rect 790 14374 833 14438
rect 1150 14437 1216 14438
rect 725 14373 791 14374
rect 1108 14373 1151 14437
rect 1215 14373 1258 14437
rect 1751 14386 1794 14449
rect 1788 14385 1794 14386
rect 1858 14386 1901 14449
rect 2999 14449 3149 14450
rect 2999 14386 3042 14449
rect 1858 14385 1864 14386
rect 3036 14385 3042 14386
rect 3106 14386 3149 14449
rect 3106 14385 3112 14386
rect 1793 14384 1859 14385
rect 3041 14384 3107 14385
rect 1150 14372 1216 14373
rect 1150 14067 1216 14068
rect 725 14066 791 14067
rect 683 14002 726 14066
rect 790 14002 833 14066
rect 1108 14003 1151 14067
rect 1215 14003 1258 14067
rect 1793 14055 1859 14056
rect 3041 14055 3107 14056
rect 1788 14054 1794 14055
rect 1150 14002 1216 14003
rect 725 14001 791 14002
rect 1751 13991 1794 14054
rect 1858 14054 1864 14055
rect 3036 14054 3042 14055
rect 1858 13991 1901 14054
rect 1751 13990 1901 13991
rect 2999 13991 3042 14054
rect 3106 14054 3112 14055
rect 3106 13991 3149 14054
rect 2999 13990 3149 13991
rect 1751 13659 1901 13660
rect 725 13648 791 13649
rect 683 13584 726 13648
rect 790 13584 833 13648
rect 1150 13647 1216 13648
rect 725 13583 791 13584
rect 1108 13583 1151 13647
rect 1215 13583 1258 13647
rect 1751 13596 1794 13659
rect 1788 13595 1794 13596
rect 1858 13596 1901 13659
rect 2999 13659 3149 13660
rect 2999 13596 3042 13659
rect 1858 13595 1864 13596
rect 3036 13595 3042 13596
rect 3106 13596 3149 13659
rect 3106 13595 3112 13596
rect 1793 13594 1859 13595
rect 3041 13594 3107 13595
rect 1150 13582 1216 13583
rect 1150 13277 1216 13278
rect 725 13276 791 13277
rect 683 13212 726 13276
rect 790 13212 833 13276
rect 1108 13213 1151 13277
rect 1215 13213 1258 13277
rect 1793 13265 1859 13266
rect 3041 13265 3107 13266
rect 1788 13264 1794 13265
rect 1150 13212 1216 13213
rect 725 13211 791 13212
rect 1751 13201 1794 13264
rect 1858 13264 1864 13265
rect 3036 13264 3042 13265
rect 1858 13201 1901 13264
rect 1751 13200 1901 13201
rect 2999 13201 3042 13264
rect 3106 13264 3112 13265
rect 3106 13201 3149 13264
rect 2999 13200 3149 13201
rect 1751 12869 1901 12870
rect 725 12858 791 12859
rect 683 12794 726 12858
rect 790 12794 833 12858
rect 1150 12857 1216 12858
rect 725 12793 791 12794
rect 1108 12793 1151 12857
rect 1215 12793 1258 12857
rect 1751 12806 1794 12869
rect 1788 12805 1794 12806
rect 1858 12806 1901 12869
rect 2999 12869 3149 12870
rect 2999 12806 3042 12869
rect 1858 12805 1864 12806
rect 3036 12805 3042 12806
rect 3106 12806 3149 12869
rect 3106 12805 3112 12806
rect 1793 12804 1859 12805
rect 3041 12804 3107 12805
rect 1150 12792 1216 12793
rect 1150 12487 1216 12488
rect 725 12486 791 12487
rect 683 12422 726 12486
rect 790 12422 833 12486
rect 1108 12423 1151 12487
rect 1215 12423 1258 12487
rect 1793 12475 1859 12476
rect 3041 12475 3107 12476
rect 1788 12474 1794 12475
rect 1150 12422 1216 12423
rect 725 12421 791 12422
rect 1751 12411 1794 12474
rect 1858 12474 1864 12475
rect 3036 12474 3042 12475
rect 1858 12411 1901 12474
rect 1751 12410 1901 12411
rect 2999 12411 3042 12474
rect 3106 12474 3112 12475
rect 3106 12411 3149 12474
rect 2999 12410 3149 12411
rect 1751 12079 1901 12080
rect 725 12068 791 12069
rect 683 12004 726 12068
rect 790 12004 833 12068
rect 1150 12067 1216 12068
rect 725 12003 791 12004
rect 1108 12003 1151 12067
rect 1215 12003 1258 12067
rect 1751 12016 1794 12079
rect 1788 12015 1794 12016
rect 1858 12016 1901 12079
rect 2999 12079 3149 12080
rect 2999 12016 3042 12079
rect 1858 12015 1864 12016
rect 3036 12015 3042 12016
rect 3106 12016 3149 12079
rect 3106 12015 3112 12016
rect 1793 12014 1859 12015
rect 3041 12014 3107 12015
rect 1150 12002 1216 12003
rect 1150 11697 1216 11698
rect 725 11696 791 11697
rect 683 11632 726 11696
rect 790 11632 833 11696
rect 1108 11633 1151 11697
rect 1215 11633 1258 11697
rect 1793 11685 1859 11686
rect 3041 11685 3107 11686
rect 1788 11684 1794 11685
rect 1150 11632 1216 11633
rect 725 11631 791 11632
rect 1751 11621 1794 11684
rect 1858 11684 1864 11685
rect 3036 11684 3042 11685
rect 1858 11621 1901 11684
rect 1751 11620 1901 11621
rect 2999 11621 3042 11684
rect 3106 11684 3112 11685
rect 3106 11621 3149 11684
rect 2999 11620 3149 11621
rect 1751 11289 1901 11290
rect 725 11278 791 11279
rect 683 11214 726 11278
rect 790 11214 833 11278
rect 1150 11277 1216 11278
rect 725 11213 791 11214
rect 1108 11213 1151 11277
rect 1215 11213 1258 11277
rect 1751 11226 1794 11289
rect 1788 11225 1794 11226
rect 1858 11226 1901 11289
rect 2999 11289 3149 11290
rect 2999 11226 3042 11289
rect 1858 11225 1864 11226
rect 3036 11225 3042 11226
rect 3106 11226 3149 11289
rect 3106 11225 3112 11226
rect 1793 11224 1859 11225
rect 3041 11224 3107 11225
rect 1150 11212 1216 11213
rect 1150 10907 1216 10908
rect 725 10906 791 10907
rect 683 10842 726 10906
rect 790 10842 833 10906
rect 1108 10843 1151 10907
rect 1215 10843 1258 10907
rect 1793 10895 1859 10896
rect 3041 10895 3107 10896
rect 1788 10894 1794 10895
rect 1150 10842 1216 10843
rect 725 10841 791 10842
rect 1751 10831 1794 10894
rect 1858 10894 1864 10895
rect 3036 10894 3042 10895
rect 1858 10831 1901 10894
rect 1751 10830 1901 10831
rect 2999 10831 3042 10894
rect 3106 10894 3112 10895
rect 3106 10831 3149 10894
rect 2999 10830 3149 10831
rect 1751 10499 1901 10500
rect 725 10488 791 10489
rect 683 10424 726 10488
rect 790 10424 833 10488
rect 1150 10487 1216 10488
rect 725 10423 791 10424
rect 1108 10423 1151 10487
rect 1215 10423 1258 10487
rect 1751 10436 1794 10499
rect 1788 10435 1794 10436
rect 1858 10436 1901 10499
rect 2999 10499 3149 10500
rect 2999 10436 3042 10499
rect 1858 10435 1864 10436
rect 3036 10435 3042 10436
rect 3106 10436 3149 10499
rect 3106 10435 3112 10436
rect 1793 10434 1859 10435
rect 3041 10434 3107 10435
rect 1150 10422 1216 10423
rect 1150 10117 1216 10118
rect 725 10116 791 10117
rect 683 10052 726 10116
rect 790 10052 833 10116
rect 1108 10053 1151 10117
rect 1215 10053 1258 10117
rect 1793 10105 1859 10106
rect 3041 10105 3107 10106
rect 1788 10104 1794 10105
rect 1150 10052 1216 10053
rect 725 10051 791 10052
rect 1751 10041 1794 10104
rect 1858 10104 1864 10105
rect 3036 10104 3042 10105
rect 1858 10041 1901 10104
rect 1751 10040 1901 10041
rect 2999 10041 3042 10104
rect 3106 10104 3112 10105
rect 3106 10041 3149 10104
rect 2999 10040 3149 10041
rect 1751 9709 1901 9710
rect 725 9698 791 9699
rect 683 9634 726 9698
rect 790 9634 833 9698
rect 1150 9697 1216 9698
rect 725 9633 791 9634
rect 1108 9633 1151 9697
rect 1215 9633 1258 9697
rect 1751 9646 1794 9709
rect 1788 9645 1794 9646
rect 1858 9646 1901 9709
rect 2999 9709 3149 9710
rect 2999 9646 3042 9709
rect 1858 9645 1864 9646
rect 3036 9645 3042 9646
rect 3106 9646 3149 9709
rect 3106 9645 3112 9646
rect 1793 9644 1859 9645
rect 3041 9644 3107 9645
rect 1150 9632 1216 9633
rect 1150 9327 1216 9328
rect 725 9326 791 9327
rect 683 9262 726 9326
rect 790 9262 833 9326
rect 1108 9263 1151 9327
rect 1215 9263 1258 9327
rect 1793 9315 1859 9316
rect 3041 9315 3107 9316
rect 1788 9314 1794 9315
rect 1150 9262 1216 9263
rect 725 9261 791 9262
rect 1751 9251 1794 9314
rect 1858 9314 1864 9315
rect 3036 9314 3042 9315
rect 1858 9251 1901 9314
rect 1751 9250 1901 9251
rect 2999 9251 3042 9314
rect 3106 9314 3112 9315
rect 3106 9251 3149 9314
rect 2999 9250 3149 9251
rect 1751 8919 1901 8920
rect 725 8908 791 8909
rect 683 8844 726 8908
rect 790 8844 833 8908
rect 1150 8907 1216 8908
rect 725 8843 791 8844
rect 1108 8843 1151 8907
rect 1215 8843 1258 8907
rect 1751 8856 1794 8919
rect 1788 8855 1794 8856
rect 1858 8856 1901 8919
rect 2999 8919 3149 8920
rect 2999 8856 3042 8919
rect 1858 8855 1864 8856
rect 3036 8855 3042 8856
rect 3106 8856 3149 8919
rect 3106 8855 3112 8856
rect 1793 8854 1859 8855
rect 3041 8854 3107 8855
rect 1150 8842 1216 8843
rect 1150 8537 1216 8538
rect 725 8536 791 8537
rect 683 8472 726 8536
rect 790 8472 833 8536
rect 1108 8473 1151 8537
rect 1215 8473 1258 8537
rect 1793 8525 1859 8526
rect 3041 8525 3107 8526
rect 1788 8524 1794 8525
rect 1150 8472 1216 8473
rect 725 8471 791 8472
rect 1751 8461 1794 8524
rect 1858 8524 1864 8525
rect 3036 8524 3042 8525
rect 1858 8461 1901 8524
rect 1751 8460 1901 8461
rect 2999 8461 3042 8524
rect 3106 8524 3112 8525
rect 3106 8461 3149 8524
rect 2999 8460 3149 8461
rect 1751 8129 1901 8130
rect 725 8118 791 8119
rect 683 8054 726 8118
rect 790 8054 833 8118
rect 1150 8117 1216 8118
rect 725 8053 791 8054
rect 1108 8053 1151 8117
rect 1215 8053 1258 8117
rect 1751 8066 1794 8129
rect 1788 8065 1794 8066
rect 1858 8066 1901 8129
rect 2999 8129 3149 8130
rect 2999 8066 3042 8129
rect 1858 8065 1864 8066
rect 3036 8065 3042 8066
rect 3106 8066 3149 8129
rect 3106 8065 3112 8066
rect 1793 8064 1859 8065
rect 3041 8064 3107 8065
rect 1150 8052 1216 8053
rect 1150 7747 1216 7748
rect 725 7746 791 7747
rect 683 7682 726 7746
rect 790 7682 833 7746
rect 1108 7683 1151 7747
rect 1215 7683 1258 7747
rect 1793 7735 1859 7736
rect 3041 7735 3107 7736
rect 1788 7734 1794 7735
rect 1150 7682 1216 7683
rect 725 7681 791 7682
rect 1751 7671 1794 7734
rect 1858 7734 1864 7735
rect 3036 7734 3042 7735
rect 1858 7671 1901 7734
rect 1751 7670 1901 7671
rect 2999 7671 3042 7734
rect 3106 7734 3112 7735
rect 3106 7671 3149 7734
rect 2999 7670 3149 7671
rect 1751 7339 1901 7340
rect 725 7328 791 7329
rect 683 7264 726 7328
rect 790 7264 833 7328
rect 1150 7327 1216 7328
rect 725 7263 791 7264
rect 1108 7263 1151 7327
rect 1215 7263 1258 7327
rect 1751 7276 1794 7339
rect 1788 7275 1794 7276
rect 1858 7276 1901 7339
rect 2999 7339 3149 7340
rect 2999 7276 3042 7339
rect 1858 7275 1864 7276
rect 3036 7275 3042 7276
rect 3106 7276 3149 7339
rect 3106 7275 3112 7276
rect 1793 7274 1859 7275
rect 3041 7274 3107 7275
rect 1150 7262 1216 7263
rect 1150 6957 1216 6958
rect 725 6956 791 6957
rect 683 6892 726 6956
rect 790 6892 833 6956
rect 1108 6893 1151 6957
rect 1215 6893 1258 6957
rect 1793 6945 1859 6946
rect 3041 6945 3107 6946
rect 1788 6944 1794 6945
rect 1150 6892 1216 6893
rect 725 6891 791 6892
rect 1751 6881 1794 6944
rect 1858 6944 1864 6945
rect 3036 6944 3042 6945
rect 1858 6881 1901 6944
rect 1751 6880 1901 6881
rect 2999 6881 3042 6944
rect 3106 6944 3112 6945
rect 3106 6881 3149 6944
rect 2999 6880 3149 6881
rect 1751 6549 1901 6550
rect 725 6538 791 6539
rect 683 6474 726 6538
rect 790 6474 833 6538
rect 1150 6537 1216 6538
rect 725 6473 791 6474
rect 1108 6473 1151 6537
rect 1215 6473 1258 6537
rect 1751 6486 1794 6549
rect 1788 6485 1794 6486
rect 1858 6486 1901 6549
rect 2999 6549 3149 6550
rect 2999 6486 3042 6549
rect 1858 6485 1864 6486
rect 3036 6485 3042 6486
rect 3106 6486 3149 6549
rect 3106 6485 3112 6486
rect 1793 6484 1859 6485
rect 3041 6484 3107 6485
rect 1150 6472 1216 6473
rect 1150 6167 1216 6168
rect 725 6166 791 6167
rect 683 6102 726 6166
rect 790 6102 833 6166
rect 1108 6103 1151 6167
rect 1215 6103 1258 6167
rect 1793 6155 1859 6156
rect 3041 6155 3107 6156
rect 1788 6154 1794 6155
rect 1150 6102 1216 6103
rect 725 6101 791 6102
rect 1751 6091 1794 6154
rect 1858 6154 1864 6155
rect 3036 6154 3042 6155
rect 1858 6091 1901 6154
rect 1751 6090 1901 6091
rect 2999 6091 3042 6154
rect 3106 6154 3112 6155
rect 3106 6091 3149 6154
rect 2999 6090 3149 6091
rect 1751 5759 1901 5760
rect 725 5748 791 5749
rect 683 5684 726 5748
rect 790 5684 833 5748
rect 1150 5747 1216 5748
rect 725 5683 791 5684
rect 1108 5683 1151 5747
rect 1215 5683 1258 5747
rect 1751 5696 1794 5759
rect 1788 5695 1794 5696
rect 1858 5696 1901 5759
rect 2999 5759 3149 5760
rect 2999 5696 3042 5759
rect 1858 5695 1864 5696
rect 3036 5695 3042 5696
rect 3106 5696 3149 5759
rect 3106 5695 3112 5696
rect 1793 5694 1859 5695
rect 3041 5694 3107 5695
rect 1150 5682 1216 5683
rect 1150 5377 1216 5378
rect 725 5376 791 5377
rect 683 5312 726 5376
rect 790 5312 833 5376
rect 1108 5313 1151 5377
rect 1215 5313 1258 5377
rect 1793 5365 1859 5366
rect 3041 5365 3107 5366
rect 1788 5364 1794 5365
rect 1150 5312 1216 5313
rect 725 5311 791 5312
rect 1751 5301 1794 5364
rect 1858 5364 1864 5365
rect 3036 5364 3042 5365
rect 1858 5301 1901 5364
rect 1751 5300 1901 5301
rect 2999 5301 3042 5364
rect 3106 5364 3112 5365
rect 3106 5301 3149 5364
rect 2999 5300 3149 5301
rect 1751 4969 1901 4970
rect 725 4958 791 4959
rect 683 4894 726 4958
rect 790 4894 833 4958
rect 1150 4957 1216 4958
rect 725 4893 791 4894
rect 1108 4893 1151 4957
rect 1215 4893 1258 4957
rect 1751 4906 1794 4969
rect 1788 4905 1794 4906
rect 1858 4906 1901 4969
rect 2999 4969 3149 4970
rect 2999 4906 3042 4969
rect 1858 4905 1864 4906
rect 3036 4905 3042 4906
rect 3106 4906 3149 4969
rect 3106 4905 3112 4906
rect 1793 4904 1859 4905
rect 3041 4904 3107 4905
rect 1150 4892 1216 4893
rect 1150 4587 1216 4588
rect 725 4586 791 4587
rect 683 4522 726 4586
rect 790 4522 833 4586
rect 1108 4523 1151 4587
rect 1215 4523 1258 4587
rect 1793 4575 1859 4576
rect 3041 4575 3107 4576
rect 1788 4574 1794 4575
rect 1150 4522 1216 4523
rect 725 4521 791 4522
rect 1751 4511 1794 4574
rect 1858 4574 1864 4575
rect 3036 4574 3042 4575
rect 1858 4511 1901 4574
rect 1751 4510 1901 4511
rect 2999 4511 3042 4574
rect 3106 4574 3112 4575
rect 3106 4511 3149 4574
rect 2999 4510 3149 4511
rect 1751 4179 1901 4180
rect 725 4168 791 4169
rect 683 4104 726 4168
rect 790 4104 833 4168
rect 1150 4167 1216 4168
rect 725 4103 791 4104
rect 1108 4103 1151 4167
rect 1215 4103 1258 4167
rect 1751 4116 1794 4179
rect 1788 4115 1794 4116
rect 1858 4116 1901 4179
rect 2999 4179 3149 4180
rect 2999 4116 3042 4179
rect 1858 4115 1864 4116
rect 3036 4115 3042 4116
rect 3106 4116 3149 4179
rect 3106 4115 3112 4116
rect 1793 4114 1859 4115
rect 3041 4114 3107 4115
rect 1150 4102 1216 4103
rect 1150 3797 1216 3798
rect 725 3796 791 3797
rect 683 3732 726 3796
rect 790 3732 833 3796
rect 1108 3733 1151 3797
rect 1215 3733 1258 3797
rect 1793 3785 1859 3786
rect 3041 3785 3107 3786
rect 1788 3784 1794 3785
rect 1150 3732 1216 3733
rect 725 3731 791 3732
rect 1751 3721 1794 3784
rect 1858 3784 1864 3785
rect 3036 3784 3042 3785
rect 1858 3721 1901 3784
rect 1751 3720 1901 3721
rect 2999 3721 3042 3784
rect 3106 3784 3112 3785
rect 3106 3721 3149 3784
rect 2999 3720 3149 3721
rect 1751 3389 1901 3390
rect 725 3378 791 3379
rect 683 3314 726 3378
rect 790 3314 833 3378
rect 1150 3377 1216 3378
rect 725 3313 791 3314
rect 1108 3313 1151 3377
rect 1215 3313 1258 3377
rect 1751 3326 1794 3389
rect 1788 3325 1794 3326
rect 1858 3326 1901 3389
rect 2999 3389 3149 3390
rect 2999 3326 3042 3389
rect 1858 3325 1864 3326
rect 3036 3325 3042 3326
rect 3106 3326 3149 3389
rect 3106 3325 3112 3326
rect 1793 3324 1859 3325
rect 3041 3324 3107 3325
rect 1150 3312 1216 3313
rect 1150 3007 1216 3008
rect 725 3006 791 3007
rect 683 2942 726 3006
rect 790 2942 833 3006
rect 1108 2943 1151 3007
rect 1215 2943 1258 3007
rect 1793 2995 1859 2996
rect 3041 2995 3107 2996
rect 1788 2994 1794 2995
rect 1150 2942 1216 2943
rect 725 2941 791 2942
rect 1751 2931 1794 2994
rect 1858 2994 1864 2995
rect 3036 2994 3042 2995
rect 1858 2931 1901 2994
rect 1751 2930 1901 2931
rect 2999 2931 3042 2994
rect 3106 2994 3112 2995
rect 3106 2931 3149 2994
rect 2999 2930 3149 2931
rect 1751 2599 1901 2600
rect 725 2588 791 2589
rect 683 2524 726 2588
rect 790 2524 833 2588
rect 1150 2587 1216 2588
rect 725 2523 791 2524
rect 1108 2523 1151 2587
rect 1215 2523 1258 2587
rect 1751 2536 1794 2599
rect 1788 2535 1794 2536
rect 1858 2536 1901 2599
rect 2999 2599 3149 2600
rect 2999 2536 3042 2599
rect 1858 2535 1864 2536
rect 3036 2535 3042 2536
rect 3106 2536 3149 2599
rect 3106 2535 3112 2536
rect 1793 2534 1859 2535
rect 3041 2534 3107 2535
rect 1150 2522 1216 2523
rect 1150 2217 1216 2218
rect 725 2216 791 2217
rect 683 2152 726 2216
rect 790 2152 833 2216
rect 1108 2153 1151 2217
rect 1215 2153 1258 2217
rect 1793 2205 1859 2206
rect 3041 2205 3107 2206
rect 1788 2204 1794 2205
rect 1150 2152 1216 2153
rect 725 2151 791 2152
rect 1751 2141 1794 2204
rect 1858 2204 1864 2205
rect 3036 2204 3042 2205
rect 1858 2141 1901 2204
rect 1751 2140 1901 2141
rect 2999 2141 3042 2204
rect 3106 2204 3112 2205
rect 3106 2141 3149 2204
rect 2999 2140 3149 2141
rect 1751 1809 1901 1810
rect 725 1798 791 1799
rect 683 1734 726 1798
rect 790 1734 833 1798
rect 1150 1797 1216 1798
rect 725 1733 791 1734
rect 1108 1733 1151 1797
rect 1215 1733 1258 1797
rect 1751 1746 1794 1809
rect 1788 1745 1794 1746
rect 1858 1746 1901 1809
rect 2999 1809 3149 1810
rect 2999 1746 3042 1809
rect 1858 1745 1864 1746
rect 3036 1745 3042 1746
rect 3106 1746 3149 1809
rect 3106 1745 3112 1746
rect 1793 1744 1859 1745
rect 3041 1744 3107 1745
rect 1150 1732 1216 1733
rect 1150 1427 1216 1428
rect 725 1426 791 1427
rect 683 1362 726 1426
rect 790 1362 833 1426
rect 1108 1363 1151 1427
rect 1215 1363 1258 1427
rect 1793 1415 1859 1416
rect 3041 1415 3107 1416
rect 1788 1414 1794 1415
rect 1150 1362 1216 1363
rect 725 1361 791 1362
rect 1751 1351 1794 1414
rect 1858 1414 1864 1415
rect 3036 1414 3042 1415
rect 1858 1351 1901 1414
rect 1751 1350 1901 1351
rect 2999 1351 3042 1414
rect 3106 1414 3112 1415
rect 3106 1351 3149 1414
rect 2999 1350 3149 1351
rect 1751 1019 1901 1020
rect 725 1008 791 1009
rect 683 944 726 1008
rect 790 944 833 1008
rect 1150 1007 1216 1008
rect 725 943 791 944
rect 1108 943 1151 1007
rect 1215 943 1258 1007
rect 1751 956 1794 1019
rect 1788 955 1794 956
rect 1858 956 1901 1019
rect 2999 1019 3149 1020
rect 2999 956 3042 1019
rect 1858 955 1864 956
rect 3036 955 3042 956
rect 3106 956 3149 1019
rect 3106 955 3112 956
rect 1793 954 1859 955
rect 3041 954 3107 955
rect 1150 942 1216 943
rect 1150 637 1216 638
rect 725 636 791 637
rect 683 572 726 636
rect 790 572 833 636
rect 1108 573 1151 637
rect 1215 573 1258 637
rect 1793 625 1859 626
rect 3041 625 3107 626
rect 1788 624 1794 625
rect 1150 572 1216 573
rect 725 571 791 572
rect 1751 561 1794 624
rect 1858 624 1864 625
rect 3036 624 3042 625
rect 1858 561 1901 624
rect 1751 560 1901 561
rect 2999 561 3042 624
rect 3106 624 3112 625
rect 3106 561 3149 624
rect 2999 560 3149 561
rect 1751 229 1901 230
rect 725 218 791 219
rect 683 154 726 218
rect 790 154 833 218
rect 1150 217 1216 218
rect 725 153 791 154
rect 1108 153 1151 217
rect 1215 153 1258 217
rect 1751 166 1794 229
rect 1788 165 1794 166
rect 1858 166 1901 229
rect 2999 229 3149 230
rect 2999 166 3042 229
rect 1858 165 1864 166
rect 3036 165 3042 166
rect 3106 166 3149 229
rect 3106 165 3112 166
rect 1793 164 1859 165
rect 3041 164 3107 165
rect 1150 152 1216 153
<< via3 >>
rect 726 25122 790 25126
rect 726 25066 730 25122
rect 730 25066 786 25122
rect 786 25066 790 25122
rect 726 25062 790 25066
rect 1151 25123 1215 25127
rect 1151 25067 1155 25123
rect 1155 25067 1211 25123
rect 1211 25067 1215 25123
rect 1151 25063 1215 25067
rect 1794 25111 1858 25115
rect 1794 25055 1798 25111
rect 1798 25055 1854 25111
rect 1854 25055 1858 25111
rect 1794 25051 1858 25055
rect 3042 25111 3106 25115
rect 3042 25055 3046 25111
rect 3046 25055 3102 25111
rect 3102 25055 3106 25111
rect 3042 25051 3106 25055
rect 726 24704 790 24708
rect 726 24648 730 24704
rect 730 24648 786 24704
rect 786 24648 790 24704
rect 726 24644 790 24648
rect 1151 24703 1215 24707
rect 1151 24647 1155 24703
rect 1155 24647 1211 24703
rect 1211 24647 1215 24703
rect 1151 24643 1215 24647
rect 1794 24715 1858 24719
rect 1794 24659 1798 24715
rect 1798 24659 1854 24715
rect 1854 24659 1858 24715
rect 1794 24655 1858 24659
rect 3042 24715 3106 24719
rect 3042 24659 3046 24715
rect 3046 24659 3102 24715
rect 3102 24659 3106 24715
rect 3042 24655 3106 24659
rect 726 24332 790 24336
rect 726 24276 730 24332
rect 730 24276 786 24332
rect 786 24276 790 24332
rect 726 24272 790 24276
rect 1151 24333 1215 24337
rect 1151 24277 1155 24333
rect 1155 24277 1211 24333
rect 1211 24277 1215 24333
rect 1151 24273 1215 24277
rect 1794 24321 1858 24325
rect 1794 24265 1798 24321
rect 1798 24265 1854 24321
rect 1854 24265 1858 24321
rect 1794 24261 1858 24265
rect 3042 24321 3106 24325
rect 3042 24265 3046 24321
rect 3046 24265 3102 24321
rect 3102 24265 3106 24321
rect 3042 24261 3106 24265
rect 726 23914 790 23918
rect 726 23858 730 23914
rect 730 23858 786 23914
rect 786 23858 790 23914
rect 726 23854 790 23858
rect 1151 23913 1215 23917
rect 1151 23857 1155 23913
rect 1155 23857 1211 23913
rect 1211 23857 1215 23913
rect 1151 23853 1215 23857
rect 1794 23925 1858 23929
rect 1794 23869 1798 23925
rect 1798 23869 1854 23925
rect 1854 23869 1858 23925
rect 1794 23865 1858 23869
rect 3042 23925 3106 23929
rect 3042 23869 3046 23925
rect 3046 23869 3102 23925
rect 3102 23869 3106 23925
rect 3042 23865 3106 23869
rect 726 23542 790 23546
rect 726 23486 730 23542
rect 730 23486 786 23542
rect 786 23486 790 23542
rect 726 23482 790 23486
rect 1151 23543 1215 23547
rect 1151 23487 1155 23543
rect 1155 23487 1211 23543
rect 1211 23487 1215 23543
rect 1151 23483 1215 23487
rect 1794 23531 1858 23535
rect 1794 23475 1798 23531
rect 1798 23475 1854 23531
rect 1854 23475 1858 23531
rect 1794 23471 1858 23475
rect 3042 23531 3106 23535
rect 3042 23475 3046 23531
rect 3046 23475 3102 23531
rect 3102 23475 3106 23531
rect 3042 23471 3106 23475
rect 726 23124 790 23128
rect 726 23068 730 23124
rect 730 23068 786 23124
rect 786 23068 790 23124
rect 726 23064 790 23068
rect 1151 23123 1215 23127
rect 1151 23067 1155 23123
rect 1155 23067 1211 23123
rect 1211 23067 1215 23123
rect 1151 23063 1215 23067
rect 1794 23135 1858 23139
rect 1794 23079 1798 23135
rect 1798 23079 1854 23135
rect 1854 23079 1858 23135
rect 1794 23075 1858 23079
rect 3042 23135 3106 23139
rect 3042 23079 3046 23135
rect 3046 23079 3102 23135
rect 3102 23079 3106 23135
rect 3042 23075 3106 23079
rect 726 22752 790 22756
rect 726 22696 730 22752
rect 730 22696 786 22752
rect 786 22696 790 22752
rect 726 22692 790 22696
rect 1151 22753 1215 22757
rect 1151 22697 1155 22753
rect 1155 22697 1211 22753
rect 1211 22697 1215 22753
rect 1151 22693 1215 22697
rect 1794 22741 1858 22745
rect 1794 22685 1798 22741
rect 1798 22685 1854 22741
rect 1854 22685 1858 22741
rect 1794 22681 1858 22685
rect 3042 22741 3106 22745
rect 3042 22685 3046 22741
rect 3046 22685 3102 22741
rect 3102 22685 3106 22741
rect 3042 22681 3106 22685
rect 726 22334 790 22338
rect 726 22278 730 22334
rect 730 22278 786 22334
rect 786 22278 790 22334
rect 726 22274 790 22278
rect 1151 22333 1215 22337
rect 1151 22277 1155 22333
rect 1155 22277 1211 22333
rect 1211 22277 1215 22333
rect 1151 22273 1215 22277
rect 1794 22345 1858 22349
rect 1794 22289 1798 22345
rect 1798 22289 1854 22345
rect 1854 22289 1858 22345
rect 1794 22285 1858 22289
rect 3042 22345 3106 22349
rect 3042 22289 3046 22345
rect 3046 22289 3102 22345
rect 3102 22289 3106 22345
rect 3042 22285 3106 22289
rect 726 21962 790 21966
rect 726 21906 730 21962
rect 730 21906 786 21962
rect 786 21906 790 21962
rect 726 21902 790 21906
rect 1151 21963 1215 21967
rect 1151 21907 1155 21963
rect 1155 21907 1211 21963
rect 1211 21907 1215 21963
rect 1151 21903 1215 21907
rect 1794 21951 1858 21955
rect 1794 21895 1798 21951
rect 1798 21895 1854 21951
rect 1854 21895 1858 21951
rect 1794 21891 1858 21895
rect 3042 21951 3106 21955
rect 3042 21895 3046 21951
rect 3046 21895 3102 21951
rect 3102 21895 3106 21951
rect 3042 21891 3106 21895
rect 726 21544 790 21548
rect 726 21488 730 21544
rect 730 21488 786 21544
rect 786 21488 790 21544
rect 726 21484 790 21488
rect 1151 21543 1215 21547
rect 1151 21487 1155 21543
rect 1155 21487 1211 21543
rect 1211 21487 1215 21543
rect 1151 21483 1215 21487
rect 1794 21555 1858 21559
rect 1794 21499 1798 21555
rect 1798 21499 1854 21555
rect 1854 21499 1858 21555
rect 1794 21495 1858 21499
rect 3042 21555 3106 21559
rect 3042 21499 3046 21555
rect 3046 21499 3102 21555
rect 3102 21499 3106 21555
rect 3042 21495 3106 21499
rect 726 21172 790 21176
rect 726 21116 730 21172
rect 730 21116 786 21172
rect 786 21116 790 21172
rect 726 21112 790 21116
rect 1151 21173 1215 21177
rect 1151 21117 1155 21173
rect 1155 21117 1211 21173
rect 1211 21117 1215 21173
rect 1151 21113 1215 21117
rect 1794 21161 1858 21165
rect 1794 21105 1798 21161
rect 1798 21105 1854 21161
rect 1854 21105 1858 21161
rect 1794 21101 1858 21105
rect 3042 21161 3106 21165
rect 3042 21105 3046 21161
rect 3046 21105 3102 21161
rect 3102 21105 3106 21161
rect 3042 21101 3106 21105
rect 726 20754 790 20758
rect 726 20698 730 20754
rect 730 20698 786 20754
rect 786 20698 790 20754
rect 726 20694 790 20698
rect 1151 20753 1215 20757
rect 1151 20697 1155 20753
rect 1155 20697 1211 20753
rect 1211 20697 1215 20753
rect 1151 20693 1215 20697
rect 1794 20765 1858 20769
rect 1794 20709 1798 20765
rect 1798 20709 1854 20765
rect 1854 20709 1858 20765
rect 1794 20705 1858 20709
rect 3042 20765 3106 20769
rect 3042 20709 3046 20765
rect 3046 20709 3102 20765
rect 3102 20709 3106 20765
rect 3042 20705 3106 20709
rect 726 20382 790 20386
rect 726 20326 730 20382
rect 730 20326 786 20382
rect 786 20326 790 20382
rect 726 20322 790 20326
rect 1151 20383 1215 20387
rect 1151 20327 1155 20383
rect 1155 20327 1211 20383
rect 1211 20327 1215 20383
rect 1151 20323 1215 20327
rect 1794 20371 1858 20375
rect 1794 20315 1798 20371
rect 1798 20315 1854 20371
rect 1854 20315 1858 20371
rect 1794 20311 1858 20315
rect 3042 20371 3106 20375
rect 3042 20315 3046 20371
rect 3046 20315 3102 20371
rect 3102 20315 3106 20371
rect 3042 20311 3106 20315
rect 726 19964 790 19968
rect 726 19908 730 19964
rect 730 19908 786 19964
rect 786 19908 790 19964
rect 726 19904 790 19908
rect 1151 19963 1215 19967
rect 1151 19907 1155 19963
rect 1155 19907 1211 19963
rect 1211 19907 1215 19963
rect 1151 19903 1215 19907
rect 1794 19975 1858 19979
rect 1794 19919 1798 19975
rect 1798 19919 1854 19975
rect 1854 19919 1858 19975
rect 1794 19915 1858 19919
rect 3042 19975 3106 19979
rect 3042 19919 3046 19975
rect 3046 19919 3102 19975
rect 3102 19919 3106 19975
rect 3042 19915 3106 19919
rect 726 19592 790 19596
rect 726 19536 730 19592
rect 730 19536 786 19592
rect 786 19536 790 19592
rect 726 19532 790 19536
rect 1151 19593 1215 19597
rect 1151 19537 1155 19593
rect 1155 19537 1211 19593
rect 1211 19537 1215 19593
rect 1151 19533 1215 19537
rect 1794 19581 1858 19585
rect 1794 19525 1798 19581
rect 1798 19525 1854 19581
rect 1854 19525 1858 19581
rect 1794 19521 1858 19525
rect 3042 19581 3106 19585
rect 3042 19525 3046 19581
rect 3046 19525 3102 19581
rect 3102 19525 3106 19581
rect 3042 19521 3106 19525
rect 726 19174 790 19178
rect 726 19118 730 19174
rect 730 19118 786 19174
rect 786 19118 790 19174
rect 726 19114 790 19118
rect 1151 19173 1215 19177
rect 1151 19117 1155 19173
rect 1155 19117 1211 19173
rect 1211 19117 1215 19173
rect 1151 19113 1215 19117
rect 1794 19185 1858 19189
rect 1794 19129 1798 19185
rect 1798 19129 1854 19185
rect 1854 19129 1858 19185
rect 1794 19125 1858 19129
rect 3042 19185 3106 19189
rect 3042 19129 3046 19185
rect 3046 19129 3102 19185
rect 3102 19129 3106 19185
rect 3042 19125 3106 19129
rect 726 18802 790 18806
rect 726 18746 730 18802
rect 730 18746 786 18802
rect 786 18746 790 18802
rect 726 18742 790 18746
rect 1151 18803 1215 18807
rect 1151 18747 1155 18803
rect 1155 18747 1211 18803
rect 1211 18747 1215 18803
rect 1151 18743 1215 18747
rect 1794 18791 1858 18795
rect 1794 18735 1798 18791
rect 1798 18735 1854 18791
rect 1854 18735 1858 18791
rect 1794 18731 1858 18735
rect 3042 18791 3106 18795
rect 3042 18735 3046 18791
rect 3046 18735 3102 18791
rect 3102 18735 3106 18791
rect 3042 18731 3106 18735
rect 726 18384 790 18388
rect 726 18328 730 18384
rect 730 18328 786 18384
rect 786 18328 790 18384
rect 726 18324 790 18328
rect 1151 18383 1215 18387
rect 1151 18327 1155 18383
rect 1155 18327 1211 18383
rect 1211 18327 1215 18383
rect 1151 18323 1215 18327
rect 1794 18395 1858 18399
rect 1794 18339 1798 18395
rect 1798 18339 1854 18395
rect 1854 18339 1858 18395
rect 1794 18335 1858 18339
rect 3042 18395 3106 18399
rect 3042 18339 3046 18395
rect 3046 18339 3102 18395
rect 3102 18339 3106 18395
rect 3042 18335 3106 18339
rect 726 18012 790 18016
rect 726 17956 730 18012
rect 730 17956 786 18012
rect 786 17956 790 18012
rect 726 17952 790 17956
rect 1151 18013 1215 18017
rect 1151 17957 1155 18013
rect 1155 17957 1211 18013
rect 1211 17957 1215 18013
rect 1151 17953 1215 17957
rect 1794 18001 1858 18005
rect 1794 17945 1798 18001
rect 1798 17945 1854 18001
rect 1854 17945 1858 18001
rect 1794 17941 1858 17945
rect 3042 18001 3106 18005
rect 3042 17945 3046 18001
rect 3046 17945 3102 18001
rect 3102 17945 3106 18001
rect 3042 17941 3106 17945
rect 726 17594 790 17598
rect 726 17538 730 17594
rect 730 17538 786 17594
rect 786 17538 790 17594
rect 726 17534 790 17538
rect 1151 17593 1215 17597
rect 1151 17537 1155 17593
rect 1155 17537 1211 17593
rect 1211 17537 1215 17593
rect 1151 17533 1215 17537
rect 1794 17605 1858 17609
rect 1794 17549 1798 17605
rect 1798 17549 1854 17605
rect 1854 17549 1858 17605
rect 1794 17545 1858 17549
rect 3042 17605 3106 17609
rect 3042 17549 3046 17605
rect 3046 17549 3102 17605
rect 3102 17549 3106 17605
rect 3042 17545 3106 17549
rect 726 17222 790 17226
rect 726 17166 730 17222
rect 730 17166 786 17222
rect 786 17166 790 17222
rect 726 17162 790 17166
rect 1151 17223 1215 17227
rect 1151 17167 1155 17223
rect 1155 17167 1211 17223
rect 1211 17167 1215 17223
rect 1151 17163 1215 17167
rect 1794 17211 1858 17215
rect 1794 17155 1798 17211
rect 1798 17155 1854 17211
rect 1854 17155 1858 17211
rect 1794 17151 1858 17155
rect 3042 17211 3106 17215
rect 3042 17155 3046 17211
rect 3046 17155 3102 17211
rect 3102 17155 3106 17211
rect 3042 17151 3106 17155
rect 726 16804 790 16808
rect 726 16748 730 16804
rect 730 16748 786 16804
rect 786 16748 790 16804
rect 726 16744 790 16748
rect 1151 16803 1215 16807
rect 1151 16747 1155 16803
rect 1155 16747 1211 16803
rect 1211 16747 1215 16803
rect 1151 16743 1215 16747
rect 1794 16815 1858 16819
rect 1794 16759 1798 16815
rect 1798 16759 1854 16815
rect 1854 16759 1858 16815
rect 1794 16755 1858 16759
rect 3042 16815 3106 16819
rect 3042 16759 3046 16815
rect 3046 16759 3102 16815
rect 3102 16759 3106 16815
rect 3042 16755 3106 16759
rect 726 16432 790 16436
rect 726 16376 730 16432
rect 730 16376 786 16432
rect 786 16376 790 16432
rect 726 16372 790 16376
rect 1151 16433 1215 16437
rect 1151 16377 1155 16433
rect 1155 16377 1211 16433
rect 1211 16377 1215 16433
rect 1151 16373 1215 16377
rect 1794 16421 1858 16425
rect 1794 16365 1798 16421
rect 1798 16365 1854 16421
rect 1854 16365 1858 16421
rect 1794 16361 1858 16365
rect 3042 16421 3106 16425
rect 3042 16365 3046 16421
rect 3046 16365 3102 16421
rect 3102 16365 3106 16421
rect 3042 16361 3106 16365
rect 726 16014 790 16018
rect 726 15958 730 16014
rect 730 15958 786 16014
rect 786 15958 790 16014
rect 726 15954 790 15958
rect 1151 16013 1215 16017
rect 1151 15957 1155 16013
rect 1155 15957 1211 16013
rect 1211 15957 1215 16013
rect 1151 15953 1215 15957
rect 1794 16025 1858 16029
rect 1794 15969 1798 16025
rect 1798 15969 1854 16025
rect 1854 15969 1858 16025
rect 1794 15965 1858 15969
rect 3042 16025 3106 16029
rect 3042 15969 3046 16025
rect 3046 15969 3102 16025
rect 3102 15969 3106 16025
rect 3042 15965 3106 15969
rect 726 15642 790 15646
rect 726 15586 730 15642
rect 730 15586 786 15642
rect 786 15586 790 15642
rect 726 15582 790 15586
rect 1151 15643 1215 15647
rect 1151 15587 1155 15643
rect 1155 15587 1211 15643
rect 1211 15587 1215 15643
rect 1151 15583 1215 15587
rect 1794 15631 1858 15635
rect 1794 15575 1798 15631
rect 1798 15575 1854 15631
rect 1854 15575 1858 15631
rect 1794 15571 1858 15575
rect 3042 15631 3106 15635
rect 3042 15575 3046 15631
rect 3046 15575 3102 15631
rect 3102 15575 3106 15631
rect 3042 15571 3106 15575
rect 726 15224 790 15228
rect 726 15168 730 15224
rect 730 15168 786 15224
rect 786 15168 790 15224
rect 726 15164 790 15168
rect 1151 15223 1215 15227
rect 1151 15167 1155 15223
rect 1155 15167 1211 15223
rect 1211 15167 1215 15223
rect 1151 15163 1215 15167
rect 1794 15235 1858 15239
rect 1794 15179 1798 15235
rect 1798 15179 1854 15235
rect 1854 15179 1858 15235
rect 1794 15175 1858 15179
rect 3042 15235 3106 15239
rect 3042 15179 3046 15235
rect 3046 15179 3102 15235
rect 3102 15179 3106 15235
rect 3042 15175 3106 15179
rect 726 14852 790 14856
rect 726 14796 730 14852
rect 730 14796 786 14852
rect 786 14796 790 14852
rect 726 14792 790 14796
rect 1151 14853 1215 14857
rect 1151 14797 1155 14853
rect 1155 14797 1211 14853
rect 1211 14797 1215 14853
rect 1151 14793 1215 14797
rect 1794 14841 1858 14845
rect 1794 14785 1798 14841
rect 1798 14785 1854 14841
rect 1854 14785 1858 14841
rect 1794 14781 1858 14785
rect 3042 14841 3106 14845
rect 3042 14785 3046 14841
rect 3046 14785 3102 14841
rect 3102 14785 3106 14841
rect 3042 14781 3106 14785
rect 726 14434 790 14438
rect 726 14378 730 14434
rect 730 14378 786 14434
rect 786 14378 790 14434
rect 726 14374 790 14378
rect 1151 14433 1215 14437
rect 1151 14377 1155 14433
rect 1155 14377 1211 14433
rect 1211 14377 1215 14433
rect 1151 14373 1215 14377
rect 1794 14445 1858 14449
rect 1794 14389 1798 14445
rect 1798 14389 1854 14445
rect 1854 14389 1858 14445
rect 1794 14385 1858 14389
rect 3042 14445 3106 14449
rect 3042 14389 3046 14445
rect 3046 14389 3102 14445
rect 3102 14389 3106 14445
rect 3042 14385 3106 14389
rect 726 14062 790 14066
rect 726 14006 730 14062
rect 730 14006 786 14062
rect 786 14006 790 14062
rect 726 14002 790 14006
rect 1151 14063 1215 14067
rect 1151 14007 1155 14063
rect 1155 14007 1211 14063
rect 1211 14007 1215 14063
rect 1151 14003 1215 14007
rect 1794 14051 1858 14055
rect 1794 13995 1798 14051
rect 1798 13995 1854 14051
rect 1854 13995 1858 14051
rect 1794 13991 1858 13995
rect 3042 14051 3106 14055
rect 3042 13995 3046 14051
rect 3046 13995 3102 14051
rect 3102 13995 3106 14051
rect 3042 13991 3106 13995
rect 726 13644 790 13648
rect 726 13588 730 13644
rect 730 13588 786 13644
rect 786 13588 790 13644
rect 726 13584 790 13588
rect 1151 13643 1215 13647
rect 1151 13587 1155 13643
rect 1155 13587 1211 13643
rect 1211 13587 1215 13643
rect 1151 13583 1215 13587
rect 1794 13655 1858 13659
rect 1794 13599 1798 13655
rect 1798 13599 1854 13655
rect 1854 13599 1858 13655
rect 1794 13595 1858 13599
rect 3042 13655 3106 13659
rect 3042 13599 3046 13655
rect 3046 13599 3102 13655
rect 3102 13599 3106 13655
rect 3042 13595 3106 13599
rect 726 13272 790 13276
rect 726 13216 730 13272
rect 730 13216 786 13272
rect 786 13216 790 13272
rect 726 13212 790 13216
rect 1151 13273 1215 13277
rect 1151 13217 1155 13273
rect 1155 13217 1211 13273
rect 1211 13217 1215 13273
rect 1151 13213 1215 13217
rect 1794 13261 1858 13265
rect 1794 13205 1798 13261
rect 1798 13205 1854 13261
rect 1854 13205 1858 13261
rect 1794 13201 1858 13205
rect 3042 13261 3106 13265
rect 3042 13205 3046 13261
rect 3046 13205 3102 13261
rect 3102 13205 3106 13261
rect 3042 13201 3106 13205
rect 726 12854 790 12858
rect 726 12798 730 12854
rect 730 12798 786 12854
rect 786 12798 790 12854
rect 726 12794 790 12798
rect 1151 12853 1215 12857
rect 1151 12797 1155 12853
rect 1155 12797 1211 12853
rect 1211 12797 1215 12853
rect 1151 12793 1215 12797
rect 1794 12865 1858 12869
rect 1794 12809 1798 12865
rect 1798 12809 1854 12865
rect 1854 12809 1858 12865
rect 1794 12805 1858 12809
rect 3042 12865 3106 12869
rect 3042 12809 3046 12865
rect 3046 12809 3102 12865
rect 3102 12809 3106 12865
rect 3042 12805 3106 12809
rect 726 12482 790 12486
rect 726 12426 730 12482
rect 730 12426 786 12482
rect 786 12426 790 12482
rect 726 12422 790 12426
rect 1151 12483 1215 12487
rect 1151 12427 1155 12483
rect 1155 12427 1211 12483
rect 1211 12427 1215 12483
rect 1151 12423 1215 12427
rect 1794 12471 1858 12475
rect 1794 12415 1798 12471
rect 1798 12415 1854 12471
rect 1854 12415 1858 12471
rect 1794 12411 1858 12415
rect 3042 12471 3106 12475
rect 3042 12415 3046 12471
rect 3046 12415 3102 12471
rect 3102 12415 3106 12471
rect 3042 12411 3106 12415
rect 726 12064 790 12068
rect 726 12008 730 12064
rect 730 12008 786 12064
rect 786 12008 790 12064
rect 726 12004 790 12008
rect 1151 12063 1215 12067
rect 1151 12007 1155 12063
rect 1155 12007 1211 12063
rect 1211 12007 1215 12063
rect 1151 12003 1215 12007
rect 1794 12075 1858 12079
rect 1794 12019 1798 12075
rect 1798 12019 1854 12075
rect 1854 12019 1858 12075
rect 1794 12015 1858 12019
rect 3042 12075 3106 12079
rect 3042 12019 3046 12075
rect 3046 12019 3102 12075
rect 3102 12019 3106 12075
rect 3042 12015 3106 12019
rect 726 11692 790 11696
rect 726 11636 730 11692
rect 730 11636 786 11692
rect 786 11636 790 11692
rect 726 11632 790 11636
rect 1151 11693 1215 11697
rect 1151 11637 1155 11693
rect 1155 11637 1211 11693
rect 1211 11637 1215 11693
rect 1151 11633 1215 11637
rect 1794 11681 1858 11685
rect 1794 11625 1798 11681
rect 1798 11625 1854 11681
rect 1854 11625 1858 11681
rect 1794 11621 1858 11625
rect 3042 11681 3106 11685
rect 3042 11625 3046 11681
rect 3046 11625 3102 11681
rect 3102 11625 3106 11681
rect 3042 11621 3106 11625
rect 726 11274 790 11278
rect 726 11218 730 11274
rect 730 11218 786 11274
rect 786 11218 790 11274
rect 726 11214 790 11218
rect 1151 11273 1215 11277
rect 1151 11217 1155 11273
rect 1155 11217 1211 11273
rect 1211 11217 1215 11273
rect 1151 11213 1215 11217
rect 1794 11285 1858 11289
rect 1794 11229 1798 11285
rect 1798 11229 1854 11285
rect 1854 11229 1858 11285
rect 1794 11225 1858 11229
rect 3042 11285 3106 11289
rect 3042 11229 3046 11285
rect 3046 11229 3102 11285
rect 3102 11229 3106 11285
rect 3042 11225 3106 11229
rect 726 10902 790 10906
rect 726 10846 730 10902
rect 730 10846 786 10902
rect 786 10846 790 10902
rect 726 10842 790 10846
rect 1151 10903 1215 10907
rect 1151 10847 1155 10903
rect 1155 10847 1211 10903
rect 1211 10847 1215 10903
rect 1151 10843 1215 10847
rect 1794 10891 1858 10895
rect 1794 10835 1798 10891
rect 1798 10835 1854 10891
rect 1854 10835 1858 10891
rect 1794 10831 1858 10835
rect 3042 10891 3106 10895
rect 3042 10835 3046 10891
rect 3046 10835 3102 10891
rect 3102 10835 3106 10891
rect 3042 10831 3106 10835
rect 726 10484 790 10488
rect 726 10428 730 10484
rect 730 10428 786 10484
rect 786 10428 790 10484
rect 726 10424 790 10428
rect 1151 10483 1215 10487
rect 1151 10427 1155 10483
rect 1155 10427 1211 10483
rect 1211 10427 1215 10483
rect 1151 10423 1215 10427
rect 1794 10495 1858 10499
rect 1794 10439 1798 10495
rect 1798 10439 1854 10495
rect 1854 10439 1858 10495
rect 1794 10435 1858 10439
rect 3042 10495 3106 10499
rect 3042 10439 3046 10495
rect 3046 10439 3102 10495
rect 3102 10439 3106 10495
rect 3042 10435 3106 10439
rect 726 10112 790 10116
rect 726 10056 730 10112
rect 730 10056 786 10112
rect 786 10056 790 10112
rect 726 10052 790 10056
rect 1151 10113 1215 10117
rect 1151 10057 1155 10113
rect 1155 10057 1211 10113
rect 1211 10057 1215 10113
rect 1151 10053 1215 10057
rect 1794 10101 1858 10105
rect 1794 10045 1798 10101
rect 1798 10045 1854 10101
rect 1854 10045 1858 10101
rect 1794 10041 1858 10045
rect 3042 10101 3106 10105
rect 3042 10045 3046 10101
rect 3046 10045 3102 10101
rect 3102 10045 3106 10101
rect 3042 10041 3106 10045
rect 726 9694 790 9698
rect 726 9638 730 9694
rect 730 9638 786 9694
rect 786 9638 790 9694
rect 726 9634 790 9638
rect 1151 9693 1215 9697
rect 1151 9637 1155 9693
rect 1155 9637 1211 9693
rect 1211 9637 1215 9693
rect 1151 9633 1215 9637
rect 1794 9705 1858 9709
rect 1794 9649 1798 9705
rect 1798 9649 1854 9705
rect 1854 9649 1858 9705
rect 1794 9645 1858 9649
rect 3042 9705 3106 9709
rect 3042 9649 3046 9705
rect 3046 9649 3102 9705
rect 3102 9649 3106 9705
rect 3042 9645 3106 9649
rect 726 9322 790 9326
rect 726 9266 730 9322
rect 730 9266 786 9322
rect 786 9266 790 9322
rect 726 9262 790 9266
rect 1151 9323 1215 9327
rect 1151 9267 1155 9323
rect 1155 9267 1211 9323
rect 1211 9267 1215 9323
rect 1151 9263 1215 9267
rect 1794 9311 1858 9315
rect 1794 9255 1798 9311
rect 1798 9255 1854 9311
rect 1854 9255 1858 9311
rect 1794 9251 1858 9255
rect 3042 9311 3106 9315
rect 3042 9255 3046 9311
rect 3046 9255 3102 9311
rect 3102 9255 3106 9311
rect 3042 9251 3106 9255
rect 726 8904 790 8908
rect 726 8848 730 8904
rect 730 8848 786 8904
rect 786 8848 790 8904
rect 726 8844 790 8848
rect 1151 8903 1215 8907
rect 1151 8847 1155 8903
rect 1155 8847 1211 8903
rect 1211 8847 1215 8903
rect 1151 8843 1215 8847
rect 1794 8915 1858 8919
rect 1794 8859 1798 8915
rect 1798 8859 1854 8915
rect 1854 8859 1858 8915
rect 1794 8855 1858 8859
rect 3042 8915 3106 8919
rect 3042 8859 3046 8915
rect 3046 8859 3102 8915
rect 3102 8859 3106 8915
rect 3042 8855 3106 8859
rect 726 8532 790 8536
rect 726 8476 730 8532
rect 730 8476 786 8532
rect 786 8476 790 8532
rect 726 8472 790 8476
rect 1151 8533 1215 8537
rect 1151 8477 1155 8533
rect 1155 8477 1211 8533
rect 1211 8477 1215 8533
rect 1151 8473 1215 8477
rect 1794 8521 1858 8525
rect 1794 8465 1798 8521
rect 1798 8465 1854 8521
rect 1854 8465 1858 8521
rect 1794 8461 1858 8465
rect 3042 8521 3106 8525
rect 3042 8465 3046 8521
rect 3046 8465 3102 8521
rect 3102 8465 3106 8521
rect 3042 8461 3106 8465
rect 726 8114 790 8118
rect 726 8058 730 8114
rect 730 8058 786 8114
rect 786 8058 790 8114
rect 726 8054 790 8058
rect 1151 8113 1215 8117
rect 1151 8057 1155 8113
rect 1155 8057 1211 8113
rect 1211 8057 1215 8113
rect 1151 8053 1215 8057
rect 1794 8125 1858 8129
rect 1794 8069 1798 8125
rect 1798 8069 1854 8125
rect 1854 8069 1858 8125
rect 1794 8065 1858 8069
rect 3042 8125 3106 8129
rect 3042 8069 3046 8125
rect 3046 8069 3102 8125
rect 3102 8069 3106 8125
rect 3042 8065 3106 8069
rect 726 7742 790 7746
rect 726 7686 730 7742
rect 730 7686 786 7742
rect 786 7686 790 7742
rect 726 7682 790 7686
rect 1151 7743 1215 7747
rect 1151 7687 1155 7743
rect 1155 7687 1211 7743
rect 1211 7687 1215 7743
rect 1151 7683 1215 7687
rect 1794 7731 1858 7735
rect 1794 7675 1798 7731
rect 1798 7675 1854 7731
rect 1854 7675 1858 7731
rect 1794 7671 1858 7675
rect 3042 7731 3106 7735
rect 3042 7675 3046 7731
rect 3046 7675 3102 7731
rect 3102 7675 3106 7731
rect 3042 7671 3106 7675
rect 726 7324 790 7328
rect 726 7268 730 7324
rect 730 7268 786 7324
rect 786 7268 790 7324
rect 726 7264 790 7268
rect 1151 7323 1215 7327
rect 1151 7267 1155 7323
rect 1155 7267 1211 7323
rect 1211 7267 1215 7323
rect 1151 7263 1215 7267
rect 1794 7335 1858 7339
rect 1794 7279 1798 7335
rect 1798 7279 1854 7335
rect 1854 7279 1858 7335
rect 1794 7275 1858 7279
rect 3042 7335 3106 7339
rect 3042 7279 3046 7335
rect 3046 7279 3102 7335
rect 3102 7279 3106 7335
rect 3042 7275 3106 7279
rect 726 6952 790 6956
rect 726 6896 730 6952
rect 730 6896 786 6952
rect 786 6896 790 6952
rect 726 6892 790 6896
rect 1151 6953 1215 6957
rect 1151 6897 1155 6953
rect 1155 6897 1211 6953
rect 1211 6897 1215 6953
rect 1151 6893 1215 6897
rect 1794 6941 1858 6945
rect 1794 6885 1798 6941
rect 1798 6885 1854 6941
rect 1854 6885 1858 6941
rect 1794 6881 1858 6885
rect 3042 6941 3106 6945
rect 3042 6885 3046 6941
rect 3046 6885 3102 6941
rect 3102 6885 3106 6941
rect 3042 6881 3106 6885
rect 726 6534 790 6538
rect 726 6478 730 6534
rect 730 6478 786 6534
rect 786 6478 790 6534
rect 726 6474 790 6478
rect 1151 6533 1215 6537
rect 1151 6477 1155 6533
rect 1155 6477 1211 6533
rect 1211 6477 1215 6533
rect 1151 6473 1215 6477
rect 1794 6545 1858 6549
rect 1794 6489 1798 6545
rect 1798 6489 1854 6545
rect 1854 6489 1858 6545
rect 1794 6485 1858 6489
rect 3042 6545 3106 6549
rect 3042 6489 3046 6545
rect 3046 6489 3102 6545
rect 3102 6489 3106 6545
rect 3042 6485 3106 6489
rect 726 6162 790 6166
rect 726 6106 730 6162
rect 730 6106 786 6162
rect 786 6106 790 6162
rect 726 6102 790 6106
rect 1151 6163 1215 6167
rect 1151 6107 1155 6163
rect 1155 6107 1211 6163
rect 1211 6107 1215 6163
rect 1151 6103 1215 6107
rect 1794 6151 1858 6155
rect 1794 6095 1798 6151
rect 1798 6095 1854 6151
rect 1854 6095 1858 6151
rect 1794 6091 1858 6095
rect 3042 6151 3106 6155
rect 3042 6095 3046 6151
rect 3046 6095 3102 6151
rect 3102 6095 3106 6151
rect 3042 6091 3106 6095
rect 726 5744 790 5748
rect 726 5688 730 5744
rect 730 5688 786 5744
rect 786 5688 790 5744
rect 726 5684 790 5688
rect 1151 5743 1215 5747
rect 1151 5687 1155 5743
rect 1155 5687 1211 5743
rect 1211 5687 1215 5743
rect 1151 5683 1215 5687
rect 1794 5755 1858 5759
rect 1794 5699 1798 5755
rect 1798 5699 1854 5755
rect 1854 5699 1858 5755
rect 1794 5695 1858 5699
rect 3042 5755 3106 5759
rect 3042 5699 3046 5755
rect 3046 5699 3102 5755
rect 3102 5699 3106 5755
rect 3042 5695 3106 5699
rect 726 5372 790 5376
rect 726 5316 730 5372
rect 730 5316 786 5372
rect 786 5316 790 5372
rect 726 5312 790 5316
rect 1151 5373 1215 5377
rect 1151 5317 1155 5373
rect 1155 5317 1211 5373
rect 1211 5317 1215 5373
rect 1151 5313 1215 5317
rect 1794 5361 1858 5365
rect 1794 5305 1798 5361
rect 1798 5305 1854 5361
rect 1854 5305 1858 5361
rect 1794 5301 1858 5305
rect 3042 5361 3106 5365
rect 3042 5305 3046 5361
rect 3046 5305 3102 5361
rect 3102 5305 3106 5361
rect 3042 5301 3106 5305
rect 726 4954 790 4958
rect 726 4898 730 4954
rect 730 4898 786 4954
rect 786 4898 790 4954
rect 726 4894 790 4898
rect 1151 4953 1215 4957
rect 1151 4897 1155 4953
rect 1155 4897 1211 4953
rect 1211 4897 1215 4953
rect 1151 4893 1215 4897
rect 1794 4965 1858 4969
rect 1794 4909 1798 4965
rect 1798 4909 1854 4965
rect 1854 4909 1858 4965
rect 1794 4905 1858 4909
rect 3042 4965 3106 4969
rect 3042 4909 3046 4965
rect 3046 4909 3102 4965
rect 3102 4909 3106 4965
rect 3042 4905 3106 4909
rect 726 4582 790 4586
rect 726 4526 730 4582
rect 730 4526 786 4582
rect 786 4526 790 4582
rect 726 4522 790 4526
rect 1151 4583 1215 4587
rect 1151 4527 1155 4583
rect 1155 4527 1211 4583
rect 1211 4527 1215 4583
rect 1151 4523 1215 4527
rect 1794 4571 1858 4575
rect 1794 4515 1798 4571
rect 1798 4515 1854 4571
rect 1854 4515 1858 4571
rect 1794 4511 1858 4515
rect 3042 4571 3106 4575
rect 3042 4515 3046 4571
rect 3046 4515 3102 4571
rect 3102 4515 3106 4571
rect 3042 4511 3106 4515
rect 726 4164 790 4168
rect 726 4108 730 4164
rect 730 4108 786 4164
rect 786 4108 790 4164
rect 726 4104 790 4108
rect 1151 4163 1215 4167
rect 1151 4107 1155 4163
rect 1155 4107 1211 4163
rect 1211 4107 1215 4163
rect 1151 4103 1215 4107
rect 1794 4175 1858 4179
rect 1794 4119 1798 4175
rect 1798 4119 1854 4175
rect 1854 4119 1858 4175
rect 1794 4115 1858 4119
rect 3042 4175 3106 4179
rect 3042 4119 3046 4175
rect 3046 4119 3102 4175
rect 3102 4119 3106 4175
rect 3042 4115 3106 4119
rect 726 3792 790 3796
rect 726 3736 730 3792
rect 730 3736 786 3792
rect 786 3736 790 3792
rect 726 3732 790 3736
rect 1151 3793 1215 3797
rect 1151 3737 1155 3793
rect 1155 3737 1211 3793
rect 1211 3737 1215 3793
rect 1151 3733 1215 3737
rect 1794 3781 1858 3785
rect 1794 3725 1798 3781
rect 1798 3725 1854 3781
rect 1854 3725 1858 3781
rect 1794 3721 1858 3725
rect 3042 3781 3106 3785
rect 3042 3725 3046 3781
rect 3046 3725 3102 3781
rect 3102 3725 3106 3781
rect 3042 3721 3106 3725
rect 726 3374 790 3378
rect 726 3318 730 3374
rect 730 3318 786 3374
rect 786 3318 790 3374
rect 726 3314 790 3318
rect 1151 3373 1215 3377
rect 1151 3317 1155 3373
rect 1155 3317 1211 3373
rect 1211 3317 1215 3373
rect 1151 3313 1215 3317
rect 1794 3385 1858 3389
rect 1794 3329 1798 3385
rect 1798 3329 1854 3385
rect 1854 3329 1858 3385
rect 1794 3325 1858 3329
rect 3042 3385 3106 3389
rect 3042 3329 3046 3385
rect 3046 3329 3102 3385
rect 3102 3329 3106 3385
rect 3042 3325 3106 3329
rect 726 3002 790 3006
rect 726 2946 730 3002
rect 730 2946 786 3002
rect 786 2946 790 3002
rect 726 2942 790 2946
rect 1151 3003 1215 3007
rect 1151 2947 1155 3003
rect 1155 2947 1211 3003
rect 1211 2947 1215 3003
rect 1151 2943 1215 2947
rect 1794 2991 1858 2995
rect 1794 2935 1798 2991
rect 1798 2935 1854 2991
rect 1854 2935 1858 2991
rect 1794 2931 1858 2935
rect 3042 2991 3106 2995
rect 3042 2935 3046 2991
rect 3046 2935 3102 2991
rect 3102 2935 3106 2991
rect 3042 2931 3106 2935
rect 726 2584 790 2588
rect 726 2528 730 2584
rect 730 2528 786 2584
rect 786 2528 790 2584
rect 726 2524 790 2528
rect 1151 2583 1215 2587
rect 1151 2527 1155 2583
rect 1155 2527 1211 2583
rect 1211 2527 1215 2583
rect 1151 2523 1215 2527
rect 1794 2595 1858 2599
rect 1794 2539 1798 2595
rect 1798 2539 1854 2595
rect 1854 2539 1858 2595
rect 1794 2535 1858 2539
rect 3042 2595 3106 2599
rect 3042 2539 3046 2595
rect 3046 2539 3102 2595
rect 3102 2539 3106 2595
rect 3042 2535 3106 2539
rect 726 2212 790 2216
rect 726 2156 730 2212
rect 730 2156 786 2212
rect 786 2156 790 2212
rect 726 2152 790 2156
rect 1151 2213 1215 2217
rect 1151 2157 1155 2213
rect 1155 2157 1211 2213
rect 1211 2157 1215 2213
rect 1151 2153 1215 2157
rect 1794 2201 1858 2205
rect 1794 2145 1798 2201
rect 1798 2145 1854 2201
rect 1854 2145 1858 2201
rect 1794 2141 1858 2145
rect 3042 2201 3106 2205
rect 3042 2145 3046 2201
rect 3046 2145 3102 2201
rect 3102 2145 3106 2201
rect 3042 2141 3106 2145
rect 726 1794 790 1798
rect 726 1738 730 1794
rect 730 1738 786 1794
rect 786 1738 790 1794
rect 726 1734 790 1738
rect 1151 1793 1215 1797
rect 1151 1737 1155 1793
rect 1155 1737 1211 1793
rect 1211 1737 1215 1793
rect 1151 1733 1215 1737
rect 1794 1805 1858 1809
rect 1794 1749 1798 1805
rect 1798 1749 1854 1805
rect 1854 1749 1858 1805
rect 1794 1745 1858 1749
rect 3042 1805 3106 1809
rect 3042 1749 3046 1805
rect 3046 1749 3102 1805
rect 3102 1749 3106 1805
rect 3042 1745 3106 1749
rect 726 1422 790 1426
rect 726 1366 730 1422
rect 730 1366 786 1422
rect 786 1366 790 1422
rect 726 1362 790 1366
rect 1151 1423 1215 1427
rect 1151 1367 1155 1423
rect 1155 1367 1211 1423
rect 1211 1367 1215 1423
rect 1151 1363 1215 1367
rect 1794 1411 1858 1415
rect 1794 1355 1798 1411
rect 1798 1355 1854 1411
rect 1854 1355 1858 1411
rect 1794 1351 1858 1355
rect 3042 1411 3106 1415
rect 3042 1355 3046 1411
rect 3046 1355 3102 1411
rect 3102 1355 3106 1411
rect 3042 1351 3106 1355
rect 726 1004 790 1008
rect 726 948 730 1004
rect 730 948 786 1004
rect 786 948 790 1004
rect 726 944 790 948
rect 1151 1003 1215 1007
rect 1151 947 1155 1003
rect 1155 947 1211 1003
rect 1211 947 1215 1003
rect 1151 943 1215 947
rect 1794 1015 1858 1019
rect 1794 959 1798 1015
rect 1798 959 1854 1015
rect 1854 959 1858 1015
rect 1794 955 1858 959
rect 3042 1015 3106 1019
rect 3042 959 3046 1015
rect 3046 959 3102 1015
rect 3102 959 3106 1015
rect 3042 955 3106 959
rect 726 632 790 636
rect 726 576 730 632
rect 730 576 786 632
rect 786 576 790 632
rect 726 572 790 576
rect 1151 633 1215 637
rect 1151 577 1155 633
rect 1155 577 1211 633
rect 1211 577 1215 633
rect 1151 573 1215 577
rect 1794 621 1858 625
rect 1794 565 1798 621
rect 1798 565 1854 621
rect 1854 565 1858 621
rect 1794 561 1858 565
rect 3042 621 3106 625
rect 3042 565 3046 621
rect 3046 565 3102 621
rect 3102 565 3106 621
rect 3042 561 3106 565
rect 726 214 790 218
rect 726 158 730 214
rect 730 158 786 214
rect 786 158 790 214
rect 726 154 790 158
rect 1151 213 1215 217
rect 1151 157 1155 213
rect 1155 157 1211 213
rect 1211 157 1215 213
rect 1151 153 1215 157
rect 1794 225 1858 229
rect 1794 169 1798 225
rect 1798 169 1854 225
rect 1854 169 1858 225
rect 1794 165 1858 169
rect 3042 225 3106 229
rect 3042 169 3046 225
rect 3046 169 3102 225
rect 3102 169 3106 225
rect 3042 165 3106 169
<< metal4 >>
rect 725 25126 791 25343
rect 725 25062 726 25126
rect 790 25062 791 25126
rect 725 24708 791 25062
rect 725 24644 726 24708
rect 790 24644 791 24708
rect 725 24336 791 24644
rect 725 24272 726 24336
rect 790 24272 791 24336
rect 725 23918 791 24272
rect 725 23854 726 23918
rect 790 23854 791 23918
rect 725 23546 791 23854
rect 725 23482 726 23546
rect 790 23482 791 23546
rect 725 23128 791 23482
rect 725 23064 726 23128
rect 790 23064 791 23128
rect 725 22756 791 23064
rect 725 22692 726 22756
rect 790 22692 791 22756
rect 725 22338 791 22692
rect 725 22274 726 22338
rect 790 22274 791 22338
rect 725 21966 791 22274
rect 725 21902 726 21966
rect 790 21902 791 21966
rect 725 21548 791 21902
rect 725 21484 726 21548
rect 790 21484 791 21548
rect 725 21176 791 21484
rect 725 21112 726 21176
rect 790 21112 791 21176
rect 725 20758 791 21112
rect 725 20694 726 20758
rect 790 20694 791 20758
rect 725 20386 791 20694
rect 725 20322 726 20386
rect 790 20322 791 20386
rect 725 19968 791 20322
rect 725 19904 726 19968
rect 790 19904 791 19968
rect 725 19596 791 19904
rect 725 19532 726 19596
rect 790 19532 791 19596
rect 725 19178 791 19532
rect 725 19114 726 19178
rect 790 19114 791 19178
rect 725 18806 791 19114
rect 725 18742 726 18806
rect 790 18742 791 18806
rect 725 18388 791 18742
rect 725 18324 726 18388
rect 790 18324 791 18388
rect 725 18016 791 18324
rect 725 17952 726 18016
rect 790 17952 791 18016
rect 725 17598 791 17952
rect 725 17534 726 17598
rect 790 17534 791 17598
rect 725 17226 791 17534
rect 725 17162 726 17226
rect 790 17162 791 17226
rect 725 16808 791 17162
rect 725 16744 726 16808
rect 790 16744 791 16808
rect 725 16436 791 16744
rect 725 16372 726 16436
rect 790 16372 791 16436
rect 725 16018 791 16372
rect 725 15954 726 16018
rect 790 15954 791 16018
rect 725 15646 791 15954
rect 725 15582 726 15646
rect 790 15582 791 15646
rect 725 15228 791 15582
rect 725 15164 726 15228
rect 790 15164 791 15228
rect 725 14856 791 15164
rect 725 14792 726 14856
rect 790 14792 791 14856
rect 725 14438 791 14792
rect 725 14374 726 14438
rect 790 14374 791 14438
rect 725 14066 791 14374
rect 725 14002 726 14066
rect 790 14002 791 14066
rect 725 13648 791 14002
rect 725 13584 726 13648
rect 790 13584 791 13648
rect 725 13276 791 13584
rect 725 13212 726 13276
rect 790 13212 791 13276
rect 725 12858 791 13212
rect 725 12794 726 12858
rect 790 12794 791 12858
rect 725 12486 791 12794
rect 725 12422 726 12486
rect 790 12422 791 12486
rect 725 12068 791 12422
rect 725 12004 726 12068
rect 790 12004 791 12068
rect 725 11696 791 12004
rect 725 11632 726 11696
rect 790 11632 791 11696
rect 725 11278 791 11632
rect 725 11214 726 11278
rect 790 11214 791 11278
rect 725 10906 791 11214
rect 725 10842 726 10906
rect 790 10842 791 10906
rect 725 10488 791 10842
rect 725 10424 726 10488
rect 790 10424 791 10488
rect 725 10116 791 10424
rect 725 10052 726 10116
rect 790 10052 791 10116
rect 725 9698 791 10052
rect 725 9634 726 9698
rect 790 9634 791 9698
rect 725 9326 791 9634
rect 725 9262 726 9326
rect 790 9262 791 9326
rect 725 8908 791 9262
rect 725 8844 726 8908
rect 790 8844 791 8908
rect 725 8536 791 8844
rect 725 8472 726 8536
rect 790 8472 791 8536
rect 725 8118 791 8472
rect 725 8054 726 8118
rect 790 8054 791 8118
rect 725 7746 791 8054
rect 725 7682 726 7746
rect 790 7682 791 7746
rect 725 7328 791 7682
rect 725 7264 726 7328
rect 790 7264 791 7328
rect 725 6956 791 7264
rect 725 6892 726 6956
rect 790 6892 791 6956
rect 725 6538 791 6892
rect 725 6474 726 6538
rect 790 6474 791 6538
rect 725 6166 791 6474
rect 725 6102 726 6166
rect 790 6102 791 6166
rect 725 5748 791 6102
rect 725 5684 726 5748
rect 790 5684 791 5748
rect 725 5376 791 5684
rect 725 5312 726 5376
rect 790 5312 791 5376
rect 725 4958 791 5312
rect 725 4894 726 4958
rect 790 4894 791 4958
rect 725 4586 791 4894
rect 725 4522 726 4586
rect 790 4522 791 4586
rect 725 4168 791 4522
rect 725 4104 726 4168
rect 790 4104 791 4168
rect 725 3796 791 4104
rect 725 3732 726 3796
rect 790 3732 791 3796
rect 725 3378 791 3732
rect 725 3314 726 3378
rect 790 3314 791 3378
rect 725 3006 791 3314
rect 725 2942 726 3006
rect 790 2942 791 3006
rect 725 2588 791 2942
rect 725 2524 726 2588
rect 790 2524 791 2588
rect 725 2216 791 2524
rect 725 2152 726 2216
rect 790 2152 791 2216
rect 725 1798 791 2152
rect 725 1734 726 1798
rect 790 1734 791 1798
rect 725 1426 791 1734
rect 725 1362 726 1426
rect 790 1362 791 1426
rect 725 1008 791 1362
rect 725 944 726 1008
rect 790 944 791 1008
rect 725 636 791 944
rect 725 572 726 636
rect 790 572 791 636
rect 725 218 791 572
rect 725 154 726 218
rect 790 154 791 218
rect 725 -63 791 154
rect 1150 25127 1216 25345
rect 1150 25063 1151 25127
rect 1215 25063 1216 25127
rect 1150 24707 1216 25063
rect 1150 24643 1151 24707
rect 1215 24643 1216 24707
rect 1150 24337 1216 24643
rect 1150 24273 1151 24337
rect 1215 24273 1216 24337
rect 1150 23917 1216 24273
rect 1150 23853 1151 23917
rect 1215 23853 1216 23917
rect 1150 23547 1216 23853
rect 1150 23483 1151 23547
rect 1215 23483 1216 23547
rect 1150 23127 1216 23483
rect 1150 23063 1151 23127
rect 1215 23063 1216 23127
rect 1150 22757 1216 23063
rect 1150 22693 1151 22757
rect 1215 22693 1216 22757
rect 1150 22337 1216 22693
rect 1150 22273 1151 22337
rect 1215 22273 1216 22337
rect 1150 21967 1216 22273
rect 1150 21903 1151 21967
rect 1215 21903 1216 21967
rect 1150 21547 1216 21903
rect 1150 21483 1151 21547
rect 1215 21483 1216 21547
rect 1150 21177 1216 21483
rect 1150 21113 1151 21177
rect 1215 21113 1216 21177
rect 1150 20757 1216 21113
rect 1150 20693 1151 20757
rect 1215 20693 1216 20757
rect 1150 20387 1216 20693
rect 1150 20323 1151 20387
rect 1215 20323 1216 20387
rect 1150 19967 1216 20323
rect 1150 19903 1151 19967
rect 1215 19903 1216 19967
rect 1150 19597 1216 19903
rect 1150 19533 1151 19597
rect 1215 19533 1216 19597
rect 1150 19177 1216 19533
rect 1150 19113 1151 19177
rect 1215 19113 1216 19177
rect 1150 18807 1216 19113
rect 1150 18743 1151 18807
rect 1215 18743 1216 18807
rect 1150 18387 1216 18743
rect 1150 18323 1151 18387
rect 1215 18323 1216 18387
rect 1150 18017 1216 18323
rect 1150 17953 1151 18017
rect 1215 17953 1216 18017
rect 1150 17597 1216 17953
rect 1150 17533 1151 17597
rect 1215 17533 1216 17597
rect 1150 17227 1216 17533
rect 1150 17163 1151 17227
rect 1215 17163 1216 17227
rect 1150 16807 1216 17163
rect 1150 16743 1151 16807
rect 1215 16743 1216 16807
rect 1150 16437 1216 16743
rect 1150 16373 1151 16437
rect 1215 16373 1216 16437
rect 1150 16017 1216 16373
rect 1150 15953 1151 16017
rect 1215 15953 1216 16017
rect 1150 15647 1216 15953
rect 1150 15583 1151 15647
rect 1215 15583 1216 15647
rect 1150 15227 1216 15583
rect 1150 15163 1151 15227
rect 1215 15163 1216 15227
rect 1150 14857 1216 15163
rect 1150 14793 1151 14857
rect 1215 14793 1216 14857
rect 1150 14437 1216 14793
rect 1150 14373 1151 14437
rect 1215 14373 1216 14437
rect 1150 14067 1216 14373
rect 1150 14003 1151 14067
rect 1215 14003 1216 14067
rect 1150 13647 1216 14003
rect 1150 13583 1151 13647
rect 1215 13583 1216 13647
rect 1150 13277 1216 13583
rect 1150 13213 1151 13277
rect 1215 13213 1216 13277
rect 1150 12857 1216 13213
rect 1150 12793 1151 12857
rect 1215 12793 1216 12857
rect 1150 12487 1216 12793
rect 1150 12423 1151 12487
rect 1215 12423 1216 12487
rect 1150 12067 1216 12423
rect 1150 12003 1151 12067
rect 1215 12003 1216 12067
rect 1150 11697 1216 12003
rect 1150 11633 1151 11697
rect 1215 11633 1216 11697
rect 1150 11277 1216 11633
rect 1150 11213 1151 11277
rect 1215 11213 1216 11277
rect 1150 10907 1216 11213
rect 1150 10843 1151 10907
rect 1215 10843 1216 10907
rect 1150 10487 1216 10843
rect 1150 10423 1151 10487
rect 1215 10423 1216 10487
rect 1150 10117 1216 10423
rect 1150 10053 1151 10117
rect 1215 10053 1216 10117
rect 1150 9697 1216 10053
rect 1150 9633 1151 9697
rect 1215 9633 1216 9697
rect 1150 9327 1216 9633
rect 1150 9263 1151 9327
rect 1215 9263 1216 9327
rect 1150 8907 1216 9263
rect 1150 8843 1151 8907
rect 1215 8843 1216 8907
rect 1150 8537 1216 8843
rect 1150 8473 1151 8537
rect 1215 8473 1216 8537
rect 1150 8117 1216 8473
rect 1150 8053 1151 8117
rect 1215 8053 1216 8117
rect 1150 7747 1216 8053
rect 1150 7683 1151 7747
rect 1215 7683 1216 7747
rect 1150 7327 1216 7683
rect 1150 7263 1151 7327
rect 1215 7263 1216 7327
rect 1150 6957 1216 7263
rect 1150 6893 1151 6957
rect 1215 6893 1216 6957
rect 1150 6537 1216 6893
rect 1150 6473 1151 6537
rect 1215 6473 1216 6537
rect 1150 6167 1216 6473
rect 1150 6103 1151 6167
rect 1215 6103 1216 6167
rect 1150 5747 1216 6103
rect 1150 5683 1151 5747
rect 1215 5683 1216 5747
rect 1150 5377 1216 5683
rect 1150 5313 1151 5377
rect 1215 5313 1216 5377
rect 1150 4957 1216 5313
rect 1150 4893 1151 4957
rect 1215 4893 1216 4957
rect 1150 4587 1216 4893
rect 1150 4523 1151 4587
rect 1215 4523 1216 4587
rect 1150 4167 1216 4523
rect 1150 4103 1151 4167
rect 1215 4103 1216 4167
rect 1150 3797 1216 4103
rect 1150 3733 1151 3797
rect 1215 3733 1216 3797
rect 1150 3377 1216 3733
rect 1150 3313 1151 3377
rect 1215 3313 1216 3377
rect 1150 3007 1216 3313
rect 1150 2943 1151 3007
rect 1215 2943 1216 3007
rect 1150 2587 1216 2943
rect 1150 2523 1151 2587
rect 1215 2523 1216 2587
rect 1150 2217 1216 2523
rect 1150 2153 1151 2217
rect 1215 2153 1216 2217
rect 1150 1797 1216 2153
rect 1150 1733 1151 1797
rect 1215 1733 1216 1797
rect 1150 1427 1216 1733
rect 1150 1363 1151 1427
rect 1215 1363 1216 1427
rect 1150 1007 1216 1363
rect 1150 943 1151 1007
rect 1215 943 1216 1007
rect 1150 637 1216 943
rect 1150 573 1151 637
rect 1215 573 1216 637
rect 1150 217 1216 573
rect 1150 153 1151 217
rect 1215 153 1216 217
rect 1150 -65 1216 153
rect 1793 25115 1859 25313
rect 1793 25051 1794 25115
rect 1858 25051 1859 25115
rect 1793 24719 1859 25051
rect 1793 24655 1794 24719
rect 1858 24655 1859 24719
rect 1793 24325 1859 24655
rect 1793 24261 1794 24325
rect 1858 24261 1859 24325
rect 1793 23929 1859 24261
rect 1793 23865 1794 23929
rect 1858 23865 1859 23929
rect 1793 23535 1859 23865
rect 1793 23471 1794 23535
rect 1858 23471 1859 23535
rect 1793 23139 1859 23471
rect 1793 23075 1794 23139
rect 1858 23075 1859 23139
rect 1793 22745 1859 23075
rect 1793 22681 1794 22745
rect 1858 22681 1859 22745
rect 1793 22349 1859 22681
rect 1793 22285 1794 22349
rect 1858 22285 1859 22349
rect 1793 21955 1859 22285
rect 1793 21891 1794 21955
rect 1858 21891 1859 21955
rect 1793 21559 1859 21891
rect 1793 21495 1794 21559
rect 1858 21495 1859 21559
rect 1793 21165 1859 21495
rect 1793 21101 1794 21165
rect 1858 21101 1859 21165
rect 1793 20769 1859 21101
rect 1793 20705 1794 20769
rect 1858 20705 1859 20769
rect 1793 20375 1859 20705
rect 1793 20311 1794 20375
rect 1858 20311 1859 20375
rect 1793 19979 1859 20311
rect 1793 19915 1794 19979
rect 1858 19915 1859 19979
rect 1793 19585 1859 19915
rect 1793 19521 1794 19585
rect 1858 19521 1859 19585
rect 1793 19189 1859 19521
rect 1793 19125 1794 19189
rect 1858 19125 1859 19189
rect 1793 18795 1859 19125
rect 1793 18731 1794 18795
rect 1858 18731 1859 18795
rect 1793 18399 1859 18731
rect 1793 18335 1794 18399
rect 1858 18335 1859 18399
rect 1793 18005 1859 18335
rect 1793 17941 1794 18005
rect 1858 17941 1859 18005
rect 1793 17609 1859 17941
rect 1793 17545 1794 17609
rect 1858 17545 1859 17609
rect 1793 17215 1859 17545
rect 1793 17151 1794 17215
rect 1858 17151 1859 17215
rect 1793 16819 1859 17151
rect 1793 16755 1794 16819
rect 1858 16755 1859 16819
rect 1793 16425 1859 16755
rect 1793 16361 1794 16425
rect 1858 16361 1859 16425
rect 1793 16029 1859 16361
rect 1793 15965 1794 16029
rect 1858 15965 1859 16029
rect 1793 15635 1859 15965
rect 1793 15571 1794 15635
rect 1858 15571 1859 15635
rect 1793 15239 1859 15571
rect 1793 15175 1794 15239
rect 1858 15175 1859 15239
rect 1793 14845 1859 15175
rect 1793 14781 1794 14845
rect 1858 14781 1859 14845
rect 1793 14449 1859 14781
rect 1793 14385 1794 14449
rect 1858 14385 1859 14449
rect 1793 14055 1859 14385
rect 1793 13991 1794 14055
rect 1858 13991 1859 14055
rect 1793 13659 1859 13991
rect 1793 13595 1794 13659
rect 1858 13595 1859 13659
rect 1793 13265 1859 13595
rect 1793 13201 1794 13265
rect 1858 13201 1859 13265
rect 1793 12869 1859 13201
rect 1793 12805 1794 12869
rect 1858 12805 1859 12869
rect 1793 12475 1859 12805
rect 1793 12411 1794 12475
rect 1858 12411 1859 12475
rect 1793 12079 1859 12411
rect 1793 12015 1794 12079
rect 1858 12015 1859 12079
rect 1793 11685 1859 12015
rect 1793 11621 1794 11685
rect 1858 11621 1859 11685
rect 1793 11289 1859 11621
rect 1793 11225 1794 11289
rect 1858 11225 1859 11289
rect 1793 10895 1859 11225
rect 1793 10831 1794 10895
rect 1858 10831 1859 10895
rect 1793 10499 1859 10831
rect 1793 10435 1794 10499
rect 1858 10435 1859 10499
rect 1793 10105 1859 10435
rect 1793 10041 1794 10105
rect 1858 10041 1859 10105
rect 1793 9709 1859 10041
rect 1793 9645 1794 9709
rect 1858 9645 1859 9709
rect 1793 9315 1859 9645
rect 1793 9251 1794 9315
rect 1858 9251 1859 9315
rect 1793 8919 1859 9251
rect 1793 8855 1794 8919
rect 1858 8855 1859 8919
rect 1793 8525 1859 8855
rect 1793 8461 1794 8525
rect 1858 8461 1859 8525
rect 1793 8129 1859 8461
rect 1793 8065 1794 8129
rect 1858 8065 1859 8129
rect 1793 7735 1859 8065
rect 1793 7671 1794 7735
rect 1858 7671 1859 7735
rect 1793 7339 1859 7671
rect 1793 7275 1794 7339
rect 1858 7275 1859 7339
rect 1793 6945 1859 7275
rect 1793 6881 1794 6945
rect 1858 6881 1859 6945
rect 1793 6549 1859 6881
rect 1793 6485 1794 6549
rect 1858 6485 1859 6549
rect 1793 6155 1859 6485
rect 1793 6091 1794 6155
rect 1858 6091 1859 6155
rect 1793 5759 1859 6091
rect 1793 5695 1794 5759
rect 1858 5695 1859 5759
rect 1793 5365 1859 5695
rect 1793 5301 1794 5365
rect 1858 5301 1859 5365
rect 1793 4969 1859 5301
rect 1793 4905 1794 4969
rect 1858 4905 1859 4969
rect 1793 4575 1859 4905
rect 1793 4511 1794 4575
rect 1858 4511 1859 4575
rect 1793 4179 1859 4511
rect 1793 4115 1794 4179
rect 1858 4115 1859 4179
rect 1793 3785 1859 4115
rect 1793 3721 1794 3785
rect 1858 3721 1859 3785
rect 1793 3389 1859 3721
rect 1793 3325 1794 3389
rect 1858 3325 1859 3389
rect 1793 2995 1859 3325
rect 1793 2931 1794 2995
rect 1858 2931 1859 2995
rect 1793 2599 1859 2931
rect 1793 2535 1794 2599
rect 1858 2535 1859 2599
rect 1793 2205 1859 2535
rect 1793 2141 1794 2205
rect 1858 2141 1859 2205
rect 1793 1809 1859 2141
rect 1793 1745 1794 1809
rect 1858 1745 1859 1809
rect 1793 1415 1859 1745
rect 1793 1351 1794 1415
rect 1858 1351 1859 1415
rect 1793 1019 1859 1351
rect 1793 955 1794 1019
rect 1858 955 1859 1019
rect 1793 625 1859 955
rect 1793 561 1794 625
rect 1858 561 1859 625
rect 1793 229 1859 561
rect 1793 165 1794 229
rect 1858 165 1859 229
rect 1793 -33 1859 165
rect 3041 25115 3107 25313
rect 3041 25051 3042 25115
rect 3106 25051 3107 25115
rect 3041 24719 3107 25051
rect 3041 24655 3042 24719
rect 3106 24655 3107 24719
rect 3041 24325 3107 24655
rect 3041 24261 3042 24325
rect 3106 24261 3107 24325
rect 3041 23929 3107 24261
rect 3041 23865 3042 23929
rect 3106 23865 3107 23929
rect 3041 23535 3107 23865
rect 3041 23471 3042 23535
rect 3106 23471 3107 23535
rect 3041 23139 3107 23471
rect 3041 23075 3042 23139
rect 3106 23075 3107 23139
rect 3041 22745 3107 23075
rect 3041 22681 3042 22745
rect 3106 22681 3107 22745
rect 3041 22349 3107 22681
rect 3041 22285 3042 22349
rect 3106 22285 3107 22349
rect 3041 21955 3107 22285
rect 3041 21891 3042 21955
rect 3106 21891 3107 21955
rect 3041 21559 3107 21891
rect 3041 21495 3042 21559
rect 3106 21495 3107 21559
rect 3041 21165 3107 21495
rect 3041 21101 3042 21165
rect 3106 21101 3107 21165
rect 3041 20769 3107 21101
rect 3041 20705 3042 20769
rect 3106 20705 3107 20769
rect 3041 20375 3107 20705
rect 3041 20311 3042 20375
rect 3106 20311 3107 20375
rect 3041 19979 3107 20311
rect 3041 19915 3042 19979
rect 3106 19915 3107 19979
rect 3041 19585 3107 19915
rect 3041 19521 3042 19585
rect 3106 19521 3107 19585
rect 3041 19189 3107 19521
rect 3041 19125 3042 19189
rect 3106 19125 3107 19189
rect 3041 18795 3107 19125
rect 3041 18731 3042 18795
rect 3106 18731 3107 18795
rect 3041 18399 3107 18731
rect 3041 18335 3042 18399
rect 3106 18335 3107 18399
rect 3041 18005 3107 18335
rect 3041 17941 3042 18005
rect 3106 17941 3107 18005
rect 3041 17609 3107 17941
rect 3041 17545 3042 17609
rect 3106 17545 3107 17609
rect 3041 17215 3107 17545
rect 3041 17151 3042 17215
rect 3106 17151 3107 17215
rect 3041 16819 3107 17151
rect 3041 16755 3042 16819
rect 3106 16755 3107 16819
rect 3041 16425 3107 16755
rect 3041 16361 3042 16425
rect 3106 16361 3107 16425
rect 3041 16029 3107 16361
rect 3041 15965 3042 16029
rect 3106 15965 3107 16029
rect 3041 15635 3107 15965
rect 3041 15571 3042 15635
rect 3106 15571 3107 15635
rect 3041 15239 3107 15571
rect 3041 15175 3042 15239
rect 3106 15175 3107 15239
rect 3041 14845 3107 15175
rect 3041 14781 3042 14845
rect 3106 14781 3107 14845
rect 3041 14449 3107 14781
rect 3041 14385 3042 14449
rect 3106 14385 3107 14449
rect 3041 14055 3107 14385
rect 3041 13991 3042 14055
rect 3106 13991 3107 14055
rect 3041 13659 3107 13991
rect 3041 13595 3042 13659
rect 3106 13595 3107 13659
rect 3041 13265 3107 13595
rect 3041 13201 3042 13265
rect 3106 13201 3107 13265
rect 3041 12869 3107 13201
rect 3041 12805 3042 12869
rect 3106 12805 3107 12869
rect 3041 12475 3107 12805
rect 3041 12411 3042 12475
rect 3106 12411 3107 12475
rect 3041 12079 3107 12411
rect 3041 12015 3042 12079
rect 3106 12015 3107 12079
rect 3041 11685 3107 12015
rect 3041 11621 3042 11685
rect 3106 11621 3107 11685
rect 3041 11289 3107 11621
rect 3041 11225 3042 11289
rect 3106 11225 3107 11289
rect 3041 10895 3107 11225
rect 3041 10831 3042 10895
rect 3106 10831 3107 10895
rect 3041 10499 3107 10831
rect 3041 10435 3042 10499
rect 3106 10435 3107 10499
rect 3041 10105 3107 10435
rect 3041 10041 3042 10105
rect 3106 10041 3107 10105
rect 3041 9709 3107 10041
rect 3041 9645 3042 9709
rect 3106 9645 3107 9709
rect 3041 9315 3107 9645
rect 3041 9251 3042 9315
rect 3106 9251 3107 9315
rect 3041 8919 3107 9251
rect 3041 8855 3042 8919
rect 3106 8855 3107 8919
rect 3041 8525 3107 8855
rect 3041 8461 3042 8525
rect 3106 8461 3107 8525
rect 3041 8129 3107 8461
rect 3041 8065 3042 8129
rect 3106 8065 3107 8129
rect 3041 7735 3107 8065
rect 3041 7671 3042 7735
rect 3106 7671 3107 7735
rect 3041 7339 3107 7671
rect 3041 7275 3042 7339
rect 3106 7275 3107 7339
rect 3041 6945 3107 7275
rect 3041 6881 3042 6945
rect 3106 6881 3107 6945
rect 3041 6549 3107 6881
rect 3041 6485 3042 6549
rect 3106 6485 3107 6549
rect 3041 6155 3107 6485
rect 3041 6091 3042 6155
rect 3106 6091 3107 6155
rect 3041 5759 3107 6091
rect 3041 5695 3042 5759
rect 3106 5695 3107 5759
rect 3041 5365 3107 5695
rect 3041 5301 3042 5365
rect 3106 5301 3107 5365
rect 3041 4969 3107 5301
rect 3041 4905 3042 4969
rect 3106 4905 3107 4969
rect 3041 4575 3107 4905
rect 3041 4511 3042 4575
rect 3106 4511 3107 4575
rect 3041 4179 3107 4511
rect 3041 4115 3042 4179
rect 3106 4115 3107 4179
rect 3041 3785 3107 4115
rect 3041 3721 3042 3785
rect 3106 3721 3107 3785
rect 3041 3389 3107 3721
rect 3041 3325 3042 3389
rect 3106 3325 3107 3389
rect 3041 2995 3107 3325
rect 3041 2931 3042 2995
rect 3106 2931 3107 2995
rect 3041 2599 3107 2931
rect 3041 2535 3042 2599
rect 3106 2535 3107 2599
rect 3041 2205 3107 2535
rect 3041 2141 3042 2205
rect 3106 2141 3107 2205
rect 3041 1809 3107 2141
rect 3041 1745 3042 1809
rect 3106 1745 3107 1809
rect 3041 1415 3107 1745
rect 3041 1351 3042 1415
rect 3106 1351 3107 1415
rect 3041 1019 3107 1351
rect 3041 955 3042 1019
rect 3106 955 3107 1019
rect 3041 625 3107 955
rect 3041 561 3042 625
rect 3106 561 3107 625
rect 3041 229 3107 561
rect 3041 165 3042 229
rect 3106 165 3107 229
rect 3041 -33 3107 165
use subbyte2_wordline_driver  subbyte2_wordline_driver_0
timestamp 1543373570
transform 1 0 488 0 -1 25280
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_1
timestamp 1543373570
transform 1 0 488 0 1 24490
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_2
timestamp 1543373570
transform 1 0 488 0 -1 24490
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_3
timestamp 1543373570
transform 1 0 488 0 1 23700
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_4
timestamp 1543373570
transform 1 0 488 0 -1 23700
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_5
timestamp 1543373570
transform 1 0 488 0 1 22910
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_6
timestamp 1543373570
transform 1 0 488 0 -1 22910
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_7
timestamp 1543373570
transform 1 0 488 0 1 22120
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_8
timestamp 1543373570
transform 1 0 488 0 -1 22120
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_9
timestamp 1543373570
transform 1 0 488 0 1 21330
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_10
timestamp 1543373570
transform 1 0 488 0 -1 21330
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_11
timestamp 1543373570
transform 1 0 488 0 1 20540
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_12
timestamp 1543373570
transform 1 0 488 0 -1 20540
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_13
timestamp 1543373570
transform 1 0 488 0 1 19750
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_14
timestamp 1543373570
transform 1 0 488 0 -1 19750
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_15
timestamp 1543373570
transform 1 0 488 0 1 18960
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_16
timestamp 1543373570
transform 1 0 488 0 -1 18960
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_17
timestamp 1543373570
transform 1 0 488 0 1 18170
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_18
timestamp 1543373570
transform 1 0 488 0 -1 18170
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_19
timestamp 1543373570
transform 1 0 488 0 1 17380
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_20
timestamp 1543373570
transform 1 0 488 0 -1 17380
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_21
timestamp 1543373570
transform 1 0 488 0 1 16590
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_22
timestamp 1543373570
transform 1 0 488 0 -1 16590
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_23
timestamp 1543373570
transform 1 0 488 0 1 15800
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_24
timestamp 1543373570
transform 1 0 488 0 -1 15800
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_25
timestamp 1543373570
transform 1 0 488 0 1 15010
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_26
timestamp 1543373570
transform 1 0 488 0 -1 15010
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_27
timestamp 1543373570
transform 1 0 488 0 1 14220
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_28
timestamp 1543373570
transform 1 0 488 0 -1 14220
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_29
timestamp 1543373570
transform 1 0 488 0 1 13430
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_30
timestamp 1543373570
transform 1 0 488 0 -1 13430
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_31
timestamp 1543373570
transform 1 0 488 0 1 12640
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_32
timestamp 1543373570
transform 1 0 488 0 -1 12640
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_33
timestamp 1543373570
transform 1 0 488 0 1 11850
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_34
timestamp 1543373570
transform 1 0 488 0 -1 11850
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_35
timestamp 1543373570
transform 1 0 488 0 1 11060
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_36
timestamp 1543373570
transform 1 0 488 0 -1 11060
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_37
timestamp 1543373570
transform 1 0 488 0 1 10270
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_38
timestamp 1543373570
transform 1 0 488 0 -1 10270
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_39
timestamp 1543373570
transform 1 0 488 0 1 9480
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_40
timestamp 1543373570
transform 1 0 488 0 -1 9480
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_41
timestamp 1543373570
transform 1 0 488 0 1 8690
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_42
timestamp 1543373570
transform 1 0 488 0 -1 8690
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_43
timestamp 1543373570
transform 1 0 488 0 1 7900
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_44
timestamp 1543373570
transform 1 0 488 0 -1 7900
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_45
timestamp 1543373570
transform 1 0 488 0 1 7110
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_46
timestamp 1543373570
transform 1 0 488 0 -1 7110
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_47
timestamp 1543373570
transform 1 0 488 0 1 6320
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_48
timestamp 1543373570
transform 1 0 488 0 -1 6320
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_49
timestamp 1543373570
transform 1 0 488 0 1 5530
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_50
timestamp 1543373570
transform 1 0 488 0 -1 5530
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_51
timestamp 1543373570
transform 1 0 488 0 1 4740
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_52
timestamp 1543373570
transform 1 0 488 0 -1 4740
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_53
timestamp 1543373570
transform 1 0 488 0 1 3950
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_54
timestamp 1543373570
transform 1 0 488 0 -1 3950
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_55
timestamp 1543373570
transform 1 0 488 0 1 3160
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_56
timestamp 1543373570
transform 1 0 488 0 -1 3160
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_57
timestamp 1543373570
transform 1 0 488 0 1 2370
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_58
timestamp 1543373570
transform 1 0 488 0 -1 2370
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_59
timestamp 1543373570
transform 1 0 488 0 1 1580
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_60
timestamp 1543373570
transform 1 0 488 0 -1 1580
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_61
timestamp 1543373570
transform 1 0 488 0 1 790
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_62
timestamp 1543373570
transform 1 0 488 0 -1 790
box 70 -56 3340 490
use subbyte2_wordline_driver  subbyte2_wordline_driver_63
timestamp 1543373570
transform 1 0 488 0 1 0
box 70 -56 3340 490
<< labels >>
rlabel metal2 s 577 0 605 25280 4 en
port 3 nsew
rlabel locali s 591 299 591 299 4 in_0
port 4 nsew
rlabel locali s 3799 120 3799 120 4 wl_0
port 5 nsew
rlabel locali s 591 491 591 491 4 in_1
port 6 nsew
rlabel locali s 3799 670 3799 670 4 wl_1
port 7 nsew
rlabel locali s 591 1089 591 1089 4 in_2
port 8 nsew
rlabel locali s 3799 910 3799 910 4 wl_2
port 9 nsew
rlabel locali s 591 1281 591 1281 4 in_3
port 10 nsew
rlabel locali s 3799 1460 3799 1460 4 wl_3
port 11 nsew
rlabel locali s 591 1879 591 1879 4 in_4
port 12 nsew
rlabel locali s 3799 1700 3799 1700 4 wl_4
port 13 nsew
rlabel locali s 591 2071 591 2071 4 in_5
port 14 nsew
rlabel locali s 3799 2250 3799 2250 4 wl_5
port 15 nsew
rlabel locali s 591 2669 591 2669 4 in_6
port 16 nsew
rlabel locali s 3799 2490 3799 2490 4 wl_6
port 17 nsew
rlabel locali s 591 2861 591 2861 4 in_7
port 18 nsew
rlabel locali s 3799 3040 3799 3040 4 wl_7
port 19 nsew
rlabel locali s 591 3459 591 3459 4 in_8
port 20 nsew
rlabel locali s 3799 3280 3799 3280 4 wl_8
port 21 nsew
rlabel locali s 591 3651 591 3651 4 in_9
port 22 nsew
rlabel locali s 3799 3830 3799 3830 4 wl_9
port 23 nsew
rlabel locali s 591 4249 591 4249 4 in_10
port 24 nsew
rlabel locali s 3799 4070 3799 4070 4 wl_10
port 25 nsew
rlabel locali s 591 4441 591 4441 4 in_11
port 26 nsew
rlabel locali s 3799 4620 3799 4620 4 wl_11
port 27 nsew
rlabel locali s 591 5039 591 5039 4 in_12
port 28 nsew
rlabel locali s 3799 4860 3799 4860 4 wl_12
port 29 nsew
rlabel locali s 591 5231 591 5231 4 in_13
port 30 nsew
rlabel locali s 3799 5410 3799 5410 4 wl_13
port 31 nsew
rlabel locali s 591 5829 591 5829 4 in_14
port 32 nsew
rlabel locali s 3799 5650 3799 5650 4 wl_14
port 33 nsew
rlabel locali s 591 6021 591 6021 4 in_15
port 34 nsew
rlabel locali s 3799 6200 3799 6200 4 wl_15
port 35 nsew
rlabel locali s 591 6619 591 6619 4 in_16
port 36 nsew
rlabel locali s 3799 6440 3799 6440 4 wl_16
port 37 nsew
rlabel locali s 591 6811 591 6811 4 in_17
port 38 nsew
rlabel locali s 3799 6990 3799 6990 4 wl_17
port 39 nsew
rlabel locali s 591 7409 591 7409 4 in_18
port 40 nsew
rlabel locali s 3799 7230 3799 7230 4 wl_18
port 41 nsew
rlabel locali s 591 7601 591 7601 4 in_19
port 42 nsew
rlabel locali s 3799 7780 3799 7780 4 wl_19
port 43 nsew
rlabel locali s 591 8199 591 8199 4 in_20
port 44 nsew
rlabel locali s 3799 8020 3799 8020 4 wl_20
port 45 nsew
rlabel locali s 591 8391 591 8391 4 in_21
port 46 nsew
rlabel locali s 3799 8570 3799 8570 4 wl_21
port 47 nsew
rlabel locali s 591 8989 591 8989 4 in_22
port 48 nsew
rlabel locali s 3799 8810 3799 8810 4 wl_22
port 49 nsew
rlabel locali s 591 9181 591 9181 4 in_23
port 50 nsew
rlabel locali s 3799 9360 3799 9360 4 wl_23
port 51 nsew
rlabel locali s 591 9779 591 9779 4 in_24
port 52 nsew
rlabel locali s 3799 9600 3799 9600 4 wl_24
port 53 nsew
rlabel locali s 591 9971 591 9971 4 in_25
port 54 nsew
rlabel locali s 3799 10150 3799 10150 4 wl_25
port 55 nsew
rlabel locali s 591 10569 591 10569 4 in_26
port 56 nsew
rlabel locali s 3799 10390 3799 10390 4 wl_26
port 57 nsew
rlabel locali s 591 10761 591 10761 4 in_27
port 58 nsew
rlabel locali s 3799 10940 3799 10940 4 wl_27
port 59 nsew
rlabel locali s 591 11359 591 11359 4 in_28
port 60 nsew
rlabel locali s 3799 11180 3799 11180 4 wl_28
port 61 nsew
rlabel locali s 591 11551 591 11551 4 in_29
port 62 nsew
rlabel locali s 3799 11730 3799 11730 4 wl_29
port 63 nsew
rlabel locali s 591 12149 591 12149 4 in_30
port 64 nsew
rlabel locali s 3799 11970 3799 11970 4 wl_30
port 65 nsew
rlabel locali s 591 12341 591 12341 4 in_31
port 66 nsew
rlabel locali s 3799 12520 3799 12520 4 wl_31
port 67 nsew
rlabel locali s 591 12939 591 12939 4 in_32
port 68 nsew
rlabel locali s 3799 12760 3799 12760 4 wl_32
port 69 nsew
rlabel locali s 591 13131 591 13131 4 in_33
port 70 nsew
rlabel locali s 3799 13310 3799 13310 4 wl_33
port 71 nsew
rlabel locali s 591 13729 591 13729 4 in_34
port 72 nsew
rlabel locali s 3799 13550 3799 13550 4 wl_34
port 73 nsew
rlabel locali s 591 13921 591 13921 4 in_35
port 74 nsew
rlabel locali s 3799 14100 3799 14100 4 wl_35
port 75 nsew
rlabel locali s 591 14519 591 14519 4 in_36
port 76 nsew
rlabel locali s 3799 14340 3799 14340 4 wl_36
port 77 nsew
rlabel locali s 591 14711 591 14711 4 in_37
port 78 nsew
rlabel locali s 3799 14890 3799 14890 4 wl_37
port 79 nsew
rlabel locali s 591 15309 591 15309 4 in_38
port 80 nsew
rlabel locali s 3799 15130 3799 15130 4 wl_38
port 81 nsew
rlabel locali s 591 15501 591 15501 4 in_39
port 82 nsew
rlabel locali s 3799 15680 3799 15680 4 wl_39
port 83 nsew
rlabel locali s 591 16099 591 16099 4 in_40
port 84 nsew
rlabel locali s 3799 15920 3799 15920 4 wl_40
port 85 nsew
rlabel locali s 591 16291 591 16291 4 in_41
port 86 nsew
rlabel locali s 3799 16470 3799 16470 4 wl_41
port 87 nsew
rlabel locali s 591 16889 591 16889 4 in_42
port 88 nsew
rlabel locali s 3799 16710 3799 16710 4 wl_42
port 89 nsew
rlabel locali s 591 17081 591 17081 4 in_43
port 90 nsew
rlabel locali s 3799 17260 3799 17260 4 wl_43
port 91 nsew
rlabel locali s 591 17679 591 17679 4 in_44
port 92 nsew
rlabel locali s 3799 17500 3799 17500 4 wl_44
port 93 nsew
rlabel locali s 591 17871 591 17871 4 in_45
port 94 nsew
rlabel locali s 3799 18050 3799 18050 4 wl_45
port 95 nsew
rlabel locali s 591 18469 591 18469 4 in_46
port 96 nsew
rlabel locali s 3799 18290 3799 18290 4 wl_46
port 97 nsew
rlabel locali s 591 18661 591 18661 4 in_47
port 98 nsew
rlabel locali s 3799 18840 3799 18840 4 wl_47
port 99 nsew
rlabel locali s 591 19259 591 19259 4 in_48
port 100 nsew
rlabel locali s 3799 19080 3799 19080 4 wl_48
port 101 nsew
rlabel locali s 591 19451 591 19451 4 in_49
port 102 nsew
rlabel locali s 3799 19630 3799 19630 4 wl_49
port 103 nsew
rlabel locali s 591 20049 591 20049 4 in_50
port 104 nsew
rlabel locali s 3799 19870 3799 19870 4 wl_50
port 105 nsew
rlabel locali s 591 20241 591 20241 4 in_51
port 106 nsew
rlabel locali s 3799 20420 3799 20420 4 wl_51
port 107 nsew
rlabel locali s 591 20839 591 20839 4 in_52
port 108 nsew
rlabel locali s 3799 20660 3799 20660 4 wl_52
port 109 nsew
rlabel locali s 591 21031 591 21031 4 in_53
port 110 nsew
rlabel locali s 3799 21210 3799 21210 4 wl_53
port 111 nsew
rlabel locali s 591 21629 591 21629 4 in_54
port 112 nsew
rlabel locali s 3799 21450 3799 21450 4 wl_54
port 113 nsew
rlabel locali s 591 21821 591 21821 4 in_55
port 114 nsew
rlabel locali s 3799 22000 3799 22000 4 wl_55
port 115 nsew
rlabel locali s 591 22419 591 22419 4 in_56
port 116 nsew
rlabel locali s 3799 22240 3799 22240 4 wl_56
port 117 nsew
rlabel locali s 591 22611 591 22611 4 in_57
port 118 nsew
rlabel locali s 3799 22790 3799 22790 4 wl_57
port 119 nsew
rlabel locali s 591 23209 591 23209 4 in_58
port 120 nsew
rlabel locali s 3799 23030 3799 23030 4 wl_58
port 121 nsew
rlabel locali s 591 23401 591 23401 4 in_59
port 122 nsew
rlabel locali s 3799 23580 3799 23580 4 wl_59
port 123 nsew
rlabel locali s 591 23999 591 23999 4 in_60
port 124 nsew
rlabel locali s 3799 23820 3799 23820 4 wl_60
port 125 nsew
rlabel locali s 591 24191 591 24191 4 in_61
port 126 nsew
rlabel locali s 3799 24370 3799 24370 4 wl_61
port 127 nsew
rlabel locali s 591 24789 591 24789 4 in_62
port 128 nsew
rlabel locali s 3799 24610 3799 24610 4 wl_62
port 129 nsew
rlabel locali s 591 24981 591 24981 4 in_63
port 130 nsew
rlabel locali s 3799 25160 3799 25160 4 wl_63
port 131 nsew
rlabel metal4 s 1150 -65 1216 25345 4 vdd
port 133 nsew
rlabel metal4 s 3041 -33 3107 25313 4 vdd
port 133 nsew
rlabel metal4 s 725 -63 791 25343 4 gnd
port 135 nsew
rlabel metal4 s 1793 -33 1859 25313 4 gnd
port 135 nsew
<< properties >>
string FIXED_BBOX 0 0 3846 25280
<< end >>
