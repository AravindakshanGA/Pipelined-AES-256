magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1260 -1268 1884 1982
<< nwell >>
rect 0 0 624 722
<< scpmos >>
rect 128 416 158 526
rect 228 416 258 526
rect 128 138 158 248
<< pdiff >>
rect 68 488 128 526
rect 68 454 76 488
rect 110 454 128 488
rect 68 416 128 454
rect 158 488 228 526
rect 158 454 176 488
rect 210 454 228 488
rect 158 416 228 454
rect 258 488 318 526
rect 258 454 276 488
rect 310 454 318 488
rect 258 416 318 454
rect 68 210 128 248
rect 68 176 76 210
rect 110 176 128 210
rect 68 138 128 176
rect 158 210 218 248
rect 158 176 176 210
rect 210 176 218 210
rect 158 138 218 176
<< pdiffc >>
rect 76 454 110 488
rect 176 454 210 488
rect 276 454 310 488
rect 76 176 110 210
rect 176 176 210 210
<< nsubdiff >>
rect 168 645 218 669
rect 168 611 176 645
rect 210 611 218 645
rect 168 587 218 611
<< nsubdiffcont >>
rect 176 611 210 645
<< poly >>
rect 128 526 158 552
rect 228 526 258 552
rect 128 390 158 416
rect 228 390 258 416
rect 128 360 258 390
rect 128 248 158 360
rect 128 58 158 138
rect 125 42 191 58
rect 125 8 141 42
rect 175 8 191 42
rect 125 -8 191 8
<< polycont >>
rect 141 8 175 42
<< locali >>
rect 176 645 210 661
rect 76 488 110 504
rect 76 438 110 454
rect 176 488 210 611
rect 176 438 210 454
rect 276 488 310 504
rect 276 438 310 454
rect 76 210 110 226
rect 76 160 110 176
rect 176 210 210 226
rect 176 160 210 176
rect 141 42 175 58
rect 141 -8 175 8
<< viali >>
rect 176 611 210 645
rect 76 454 110 488
rect 276 454 310 488
rect 76 176 110 210
rect 176 176 210 210
rect 141 8 175 42
<< metal1 >>
rect 66 500 94 722
rect 164 645 222 651
rect 164 611 176 645
rect 210 611 222 645
rect 164 605 222 611
rect 530 504 558 722
rect 293 500 558 504
rect 66 488 116 500
rect 66 454 76 488
rect 110 454 116 488
rect 66 442 116 454
rect 270 488 558 500
rect 270 454 276 488
rect 310 454 558 488
rect 270 442 558 454
rect 66 222 94 442
rect 293 438 558 442
rect 530 226 558 438
rect 193 222 558 226
rect 66 210 116 222
rect 66 176 76 210
rect 110 176 116 210
rect 66 164 116 176
rect 170 210 558 222
rect 170 176 176 210
rect 210 176 558 210
rect 170 164 558 176
rect 66 0 94 164
rect 193 160 558 164
rect 126 -1 132 51
rect 184 -1 190 51
rect 530 0 558 160
<< via1 >>
rect 132 42 184 51
rect 132 8 141 42
rect 141 8 175 42
rect 175 8 184 42
rect 132 -1 184 8
<< metal2 >>
rect 132 51 184 57
rect 0 11 132 39
rect 184 11 624 39
rect 132 -7 184 -1
<< labels >>
rlabel metal2 s 0 11 624 39 4 en_bar
port 3 nsew
rlabel locali s 193 628 193 628 4 vdd
port 4 nsew
rlabel metal1 s 66 0 94 722 4 bl
port 6 nsew
rlabel metal1 s 530 0 558 722 4 br
port 8 nsew
<< properties >>
string FIXED_BBOX 105 -28 211 0
<< end >>
