magic
tech sky130A
magscale 1 2
timestamp 1714788817
<< obsli1 >>
rect 1104 2159 238832 197489
<< obsm1 >>
rect 934 1980 239094 197520
<< metal2 >>
rect 87602 199200 87658 200000
rect 88246 199200 88302 200000
rect 88890 199200 88946 200000
rect 89534 199200 89590 200000
rect 90178 199200 90234 200000
rect 90822 199200 90878 200000
rect 91466 199200 91522 200000
rect 92110 199200 92166 200000
rect 92754 199200 92810 200000
rect 93398 199200 93454 200000
rect 94042 199200 94098 200000
rect 94686 199200 94742 200000
rect 95330 199200 95386 200000
rect 95974 199200 96030 200000
rect 96618 199200 96674 200000
rect 97262 199200 97318 200000
rect 97906 199200 97962 200000
rect 98550 199200 98606 200000
rect 99194 199200 99250 200000
rect 99838 199200 99894 200000
rect 100482 199200 100538 200000
rect 101126 199200 101182 200000
rect 101770 199200 101826 200000
rect 102414 199200 102470 200000
rect 103058 199200 103114 200000
rect 103702 199200 103758 200000
rect 104346 199200 104402 200000
rect 104990 199200 105046 200000
rect 112718 199200 112774 200000
rect 113362 199200 113418 200000
rect 114006 199200 114062 200000
rect 114650 199200 114706 200000
rect 115294 199200 115350 200000
rect 115938 199200 115994 200000
rect 116582 199200 116638 200000
rect 117226 199200 117282 200000
rect 117870 199200 117926 200000
rect 118514 199200 118570 200000
rect 119158 199200 119214 200000
rect 119802 199200 119858 200000
rect 120446 199200 120502 200000
rect 121090 199200 121146 200000
rect 121734 199200 121790 200000
rect 122378 199200 122434 200000
rect 123022 199200 123078 200000
rect 123666 199200 123722 200000
rect 124310 199200 124366 200000
rect 124954 199200 125010 200000
rect 125598 199200 125654 200000
rect 126242 199200 126298 200000
rect 126886 199200 126942 200000
rect 127530 199200 127586 200000
rect 128174 199200 128230 200000
rect 128818 199200 128874 200000
rect 129462 199200 129518 200000
rect 130106 199200 130162 200000
rect 130750 199200 130806 200000
rect 131394 199200 131450 200000
rect 132038 199200 132094 200000
rect 132682 199200 132738 200000
rect 133326 199200 133382 200000
rect 133970 199200 134026 200000
rect 134614 199200 134670 200000
rect 135258 199200 135314 200000
rect 135902 199200 135958 200000
rect 136546 199200 136602 200000
rect 137190 199200 137246 200000
rect 137834 199200 137890 200000
rect 138478 199200 138534 200000
rect 139122 199200 139178 200000
rect 139766 199200 139822 200000
rect 140410 199200 140466 200000
rect 141054 199200 141110 200000
rect 141698 199200 141754 200000
rect 142342 199200 142398 200000
rect 142986 199200 143042 200000
rect 143630 199200 143686 200000
rect 144274 199200 144330 200000
rect 144918 199200 144974 200000
rect 145562 199200 145618 200000
rect 146206 199200 146262 200000
rect 146850 199200 146906 200000
rect 147494 199200 147550 200000
rect 148138 199200 148194 200000
rect 148782 199200 148838 200000
rect 149426 199200 149482 200000
rect 150070 199200 150126 200000
rect 150714 199200 150770 200000
rect 151358 199200 151414 200000
rect 152002 199200 152058 200000
rect 152646 199200 152702 200000
rect 153290 199200 153346 200000
rect 153934 199200 153990 200000
rect 154578 199200 154634 200000
rect 155222 199200 155278 200000
rect 155866 199200 155922 200000
rect 156510 199200 156566 200000
rect 157154 199200 157210 200000
rect 157798 199200 157854 200000
rect 158442 199200 158498 200000
rect 159086 199200 159142 200000
rect 159730 199200 159786 200000
rect 160374 199200 160430 200000
rect 161018 199200 161074 200000
rect 161662 199200 161718 200000
rect 162306 199200 162362 200000
rect 162950 199200 163006 200000
rect 163594 199200 163650 200000
rect 164238 199200 164294 200000
rect 164882 199200 164938 200000
rect 165526 199200 165582 200000
rect 166170 199200 166226 200000
rect 166814 199200 166870 200000
rect 167458 199200 167514 200000
rect 168102 199200 168158 200000
rect 207386 199200 207442 200000
rect 26422 0 26478 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 121090 0 121146 800
rect 121734 0 121790 800
rect 135902 0 135958 800
rect 137190 0 137246 800
<< obsm2 >>
rect 938 199144 87546 199322
rect 87714 199144 88190 199322
rect 88358 199144 88834 199322
rect 89002 199144 89478 199322
rect 89646 199144 90122 199322
rect 90290 199144 90766 199322
rect 90934 199144 91410 199322
rect 91578 199144 92054 199322
rect 92222 199144 92698 199322
rect 92866 199144 93342 199322
rect 93510 199144 93986 199322
rect 94154 199144 94630 199322
rect 94798 199144 95274 199322
rect 95442 199144 95918 199322
rect 96086 199144 96562 199322
rect 96730 199144 97206 199322
rect 97374 199144 97850 199322
rect 98018 199144 98494 199322
rect 98662 199144 99138 199322
rect 99306 199144 99782 199322
rect 99950 199144 100426 199322
rect 100594 199144 101070 199322
rect 101238 199144 101714 199322
rect 101882 199144 102358 199322
rect 102526 199144 103002 199322
rect 103170 199144 103646 199322
rect 103814 199144 104290 199322
rect 104458 199144 104934 199322
rect 105102 199144 112662 199322
rect 112830 199144 113306 199322
rect 113474 199144 113950 199322
rect 114118 199144 114594 199322
rect 114762 199144 115238 199322
rect 115406 199144 115882 199322
rect 116050 199144 116526 199322
rect 116694 199144 117170 199322
rect 117338 199144 117814 199322
rect 117982 199144 118458 199322
rect 118626 199144 119102 199322
rect 119270 199144 119746 199322
rect 119914 199144 120390 199322
rect 120558 199144 121034 199322
rect 121202 199144 121678 199322
rect 121846 199144 122322 199322
rect 122490 199144 122966 199322
rect 123134 199144 123610 199322
rect 123778 199144 124254 199322
rect 124422 199144 124898 199322
rect 125066 199144 125542 199322
rect 125710 199144 126186 199322
rect 126354 199144 126830 199322
rect 126998 199144 127474 199322
rect 127642 199144 128118 199322
rect 128286 199144 128762 199322
rect 128930 199144 129406 199322
rect 129574 199144 130050 199322
rect 130218 199144 130694 199322
rect 130862 199144 131338 199322
rect 131506 199144 131982 199322
rect 132150 199144 132626 199322
rect 132794 199144 133270 199322
rect 133438 199144 133914 199322
rect 134082 199144 134558 199322
rect 134726 199144 135202 199322
rect 135370 199144 135846 199322
rect 136014 199144 136490 199322
rect 136658 199144 137134 199322
rect 137302 199144 137778 199322
rect 137946 199144 138422 199322
rect 138590 199144 139066 199322
rect 139234 199144 139710 199322
rect 139878 199144 140354 199322
rect 140522 199144 140998 199322
rect 141166 199144 141642 199322
rect 141810 199144 142286 199322
rect 142454 199144 142930 199322
rect 143098 199144 143574 199322
rect 143742 199144 144218 199322
rect 144386 199144 144862 199322
rect 145030 199144 145506 199322
rect 145674 199144 146150 199322
rect 146318 199144 146794 199322
rect 146962 199144 147438 199322
rect 147606 199144 148082 199322
rect 148250 199144 148726 199322
rect 148894 199144 149370 199322
rect 149538 199144 150014 199322
rect 150182 199144 150658 199322
rect 150826 199144 151302 199322
rect 151470 199144 151946 199322
rect 152114 199144 152590 199322
rect 152758 199144 153234 199322
rect 153402 199144 153878 199322
rect 154046 199144 154522 199322
rect 154690 199144 155166 199322
rect 155334 199144 155810 199322
rect 155978 199144 156454 199322
rect 156622 199144 157098 199322
rect 157266 199144 157742 199322
rect 157910 199144 158386 199322
rect 158554 199144 159030 199322
rect 159198 199144 159674 199322
rect 159842 199144 160318 199322
rect 160486 199144 160962 199322
rect 161130 199144 161606 199322
rect 161774 199144 162250 199322
rect 162418 199144 162894 199322
rect 163062 199144 163538 199322
rect 163706 199144 164182 199322
rect 164350 199144 164826 199322
rect 164994 199144 165470 199322
rect 165638 199144 166114 199322
rect 166282 199144 166758 199322
rect 166926 199144 167402 199322
rect 167570 199144 168046 199322
rect 168214 199144 207330 199322
rect 207498 199144 239090 199322
rect 938 856 239090 199144
rect 938 734 26366 856
rect 26534 734 82394 856
rect 82562 734 83038 856
rect 83206 734 83682 856
rect 83850 734 84326 856
rect 84494 734 84970 856
rect 85138 734 85614 856
rect 85782 734 86258 856
rect 86426 734 86902 856
rect 87070 734 87546 856
rect 87714 734 88190 856
rect 88358 734 88834 856
rect 89002 734 89478 856
rect 89646 734 90122 856
rect 90290 734 90766 856
rect 90934 734 91410 856
rect 91578 734 92054 856
rect 92222 734 92698 856
rect 92866 734 93342 856
rect 93510 734 93986 856
rect 94154 734 94630 856
rect 94798 734 95274 856
rect 95442 734 95918 856
rect 96086 734 96562 856
rect 96730 734 97206 856
rect 97374 734 97850 856
rect 98018 734 98494 856
rect 98662 734 99138 856
rect 99306 734 99782 856
rect 99950 734 100426 856
rect 100594 734 101070 856
rect 101238 734 116526 856
rect 116694 734 117170 856
rect 117338 734 117814 856
rect 117982 734 119102 856
rect 119270 734 119746 856
rect 119914 734 120390 856
rect 120558 734 121034 856
rect 121202 734 121678 856
rect 121846 734 135846 856
rect 136014 734 137134 856
rect 137302 734 239090 856
<< metal3 >>
rect 0 138728 800 138848
rect 0 138048 800 138168
rect 0 137368 800 137488
rect 0 136688 800 136808
rect 0 114928 800 115048
rect 0 112888 800 113008
rect 239200 110168 240000 110288
rect 239200 109488 240000 109608
rect 239200 108808 240000 108928
rect 239200 108128 240000 108248
rect 239200 107448 240000 107568
rect 239200 106768 240000 106888
rect 239200 106088 240000 106208
rect 239200 105408 240000 105528
rect 239200 104728 240000 104848
rect 239200 104048 240000 104168
rect 239200 103368 240000 103488
rect 239200 102688 240000 102808
rect 239200 102008 240000 102128
rect 239200 101328 240000 101448
rect 239200 100648 240000 100768
rect 239200 99968 240000 100088
rect 0 99288 800 99408
rect 239200 99288 240000 99408
rect 0 98608 800 98728
rect 239200 98608 240000 98728
rect 239200 97928 240000 98048
rect 239200 97248 240000 97368
rect 239200 96568 240000 96688
rect 239200 95888 240000 96008
rect 239200 95208 240000 95328
rect 239200 94528 240000 94648
rect 239200 93848 240000 93968
rect 239200 93168 240000 93288
rect 239200 92488 240000 92608
rect 239200 91808 240000 91928
rect 239200 91128 240000 91248
rect 239200 90448 240000 90568
rect 239200 89768 240000 89888
rect 239200 89088 240000 89208
rect 239200 88408 240000 88528
rect 239200 87728 240000 87848
rect 239200 87048 240000 87168
rect 239200 86368 240000 86488
rect 239200 85688 240000 85808
rect 239200 85008 240000 85128
rect 239200 84328 240000 84448
rect 239200 83648 240000 83768
rect 239200 82968 240000 83088
rect 239200 82288 240000 82408
rect 239200 81608 240000 81728
rect 239200 80928 240000 81048
rect 239200 80248 240000 80368
rect 239200 79568 240000 79688
rect 239200 78888 240000 79008
rect 239200 78208 240000 78328
rect 239200 77528 240000 77648
rect 239200 76848 240000 76968
rect 239200 76168 240000 76288
rect 239200 75488 240000 75608
rect 239200 74808 240000 74928
rect 239200 74128 240000 74248
rect 239200 73448 240000 73568
rect 239200 72768 240000 72888
rect 239200 72088 240000 72208
rect 239200 71408 240000 71528
rect 239200 70728 240000 70848
rect 239200 70048 240000 70168
rect 239200 69368 240000 69488
rect 239200 68688 240000 68808
rect 239200 68008 240000 68128
rect 239200 67328 240000 67448
rect 239200 66648 240000 66768
rect 239200 65968 240000 66088
rect 239200 65288 240000 65408
rect 239200 64608 240000 64728
rect 239200 63928 240000 64048
rect 239200 63248 240000 63368
rect 239200 62568 240000 62688
rect 239200 61888 240000 62008
rect 239200 61208 240000 61328
rect 239200 60528 240000 60648
rect 239200 59848 240000 59968
rect 239200 59168 240000 59288
rect 239200 58488 240000 58608
rect 239200 57808 240000 57928
rect 239200 57128 240000 57248
rect 239200 56448 240000 56568
rect 239200 55768 240000 55888
rect 239200 55088 240000 55208
rect 239200 54408 240000 54528
rect 239200 53728 240000 53848
rect 239200 53048 240000 53168
rect 239200 52368 240000 52488
rect 239200 51688 240000 51808
rect 239200 51008 240000 51128
rect 239200 50328 240000 50448
rect 239200 49648 240000 49768
rect 239200 48968 240000 49088
rect 239200 48288 240000 48408
rect 239200 47608 240000 47728
rect 239200 46928 240000 47048
rect 239200 46248 240000 46368
rect 239200 45568 240000 45688
<< obsm3 >>
rect 798 138928 239200 197505
rect 880 138648 239200 138928
rect 798 138248 239200 138648
rect 880 137968 239200 138248
rect 798 137568 239200 137968
rect 880 137288 239200 137568
rect 798 136888 239200 137288
rect 880 136608 239200 136888
rect 798 115128 239200 136608
rect 880 114848 239200 115128
rect 798 113088 239200 114848
rect 880 112808 239200 113088
rect 798 110368 239200 112808
rect 798 110088 239120 110368
rect 798 109688 239200 110088
rect 798 109408 239120 109688
rect 798 109008 239200 109408
rect 798 108728 239120 109008
rect 798 108328 239200 108728
rect 798 108048 239120 108328
rect 798 107648 239200 108048
rect 798 107368 239120 107648
rect 798 106968 239200 107368
rect 798 106688 239120 106968
rect 798 106288 239200 106688
rect 798 106008 239120 106288
rect 798 105608 239200 106008
rect 798 105328 239120 105608
rect 798 104928 239200 105328
rect 798 104648 239120 104928
rect 798 104248 239200 104648
rect 798 103968 239120 104248
rect 798 103568 239200 103968
rect 798 103288 239120 103568
rect 798 102888 239200 103288
rect 798 102608 239120 102888
rect 798 102208 239200 102608
rect 798 101928 239120 102208
rect 798 101528 239200 101928
rect 798 101248 239120 101528
rect 798 100848 239200 101248
rect 798 100568 239120 100848
rect 798 100168 239200 100568
rect 798 99888 239120 100168
rect 798 99488 239200 99888
rect 880 99208 239120 99488
rect 798 98808 239200 99208
rect 880 98528 239120 98808
rect 798 98128 239200 98528
rect 798 97848 239120 98128
rect 798 97448 239200 97848
rect 798 97168 239120 97448
rect 798 96768 239200 97168
rect 798 96488 239120 96768
rect 798 96088 239200 96488
rect 798 95808 239120 96088
rect 798 95408 239200 95808
rect 798 95128 239120 95408
rect 798 94728 239200 95128
rect 798 94448 239120 94728
rect 798 94048 239200 94448
rect 798 93768 239120 94048
rect 798 93368 239200 93768
rect 798 93088 239120 93368
rect 798 92688 239200 93088
rect 798 92408 239120 92688
rect 798 92008 239200 92408
rect 798 91728 239120 92008
rect 798 91328 239200 91728
rect 798 91048 239120 91328
rect 798 90648 239200 91048
rect 798 90368 239120 90648
rect 798 89968 239200 90368
rect 798 89688 239120 89968
rect 798 89288 239200 89688
rect 798 89008 239120 89288
rect 798 88608 239200 89008
rect 798 88328 239120 88608
rect 798 87928 239200 88328
rect 798 87648 239120 87928
rect 798 87248 239200 87648
rect 798 86968 239120 87248
rect 798 86568 239200 86968
rect 798 86288 239120 86568
rect 798 85888 239200 86288
rect 798 85608 239120 85888
rect 798 85208 239200 85608
rect 798 84928 239120 85208
rect 798 84528 239200 84928
rect 798 84248 239120 84528
rect 798 83848 239200 84248
rect 798 83568 239120 83848
rect 798 83168 239200 83568
rect 798 82888 239120 83168
rect 798 82488 239200 82888
rect 798 82208 239120 82488
rect 798 81808 239200 82208
rect 798 81528 239120 81808
rect 798 81128 239200 81528
rect 798 80848 239120 81128
rect 798 80448 239200 80848
rect 798 80168 239120 80448
rect 798 79768 239200 80168
rect 798 79488 239120 79768
rect 798 79088 239200 79488
rect 798 78808 239120 79088
rect 798 78408 239200 78808
rect 798 78128 239120 78408
rect 798 77728 239200 78128
rect 798 77448 239120 77728
rect 798 77048 239200 77448
rect 798 76768 239120 77048
rect 798 76368 239200 76768
rect 798 76088 239120 76368
rect 798 75688 239200 76088
rect 798 75408 239120 75688
rect 798 75008 239200 75408
rect 798 74728 239120 75008
rect 798 74328 239200 74728
rect 798 74048 239120 74328
rect 798 73648 239200 74048
rect 798 73368 239120 73648
rect 798 72968 239200 73368
rect 798 72688 239120 72968
rect 798 72288 239200 72688
rect 798 72008 239120 72288
rect 798 71608 239200 72008
rect 798 71328 239120 71608
rect 798 70928 239200 71328
rect 798 70648 239120 70928
rect 798 70248 239200 70648
rect 798 69968 239120 70248
rect 798 69568 239200 69968
rect 798 69288 239120 69568
rect 798 68888 239200 69288
rect 798 68608 239120 68888
rect 798 68208 239200 68608
rect 798 67928 239120 68208
rect 798 67528 239200 67928
rect 798 67248 239120 67528
rect 798 66848 239200 67248
rect 798 66568 239120 66848
rect 798 66168 239200 66568
rect 798 65888 239120 66168
rect 798 65488 239200 65888
rect 798 65208 239120 65488
rect 798 64808 239200 65208
rect 798 64528 239120 64808
rect 798 64128 239200 64528
rect 798 63848 239120 64128
rect 798 63448 239200 63848
rect 798 63168 239120 63448
rect 798 62768 239200 63168
rect 798 62488 239120 62768
rect 798 62088 239200 62488
rect 798 61808 239120 62088
rect 798 61408 239200 61808
rect 798 61128 239120 61408
rect 798 60728 239200 61128
rect 798 60448 239120 60728
rect 798 60048 239200 60448
rect 798 59768 239120 60048
rect 798 59368 239200 59768
rect 798 59088 239120 59368
rect 798 58688 239200 59088
rect 798 58408 239120 58688
rect 798 58008 239200 58408
rect 798 57728 239120 58008
rect 798 57328 239200 57728
rect 798 57048 239120 57328
rect 798 56648 239200 57048
rect 798 56368 239120 56648
rect 798 55968 239200 56368
rect 798 55688 239120 55968
rect 798 55288 239200 55688
rect 798 55008 239120 55288
rect 798 54608 239200 55008
rect 798 54328 239120 54608
rect 798 53928 239200 54328
rect 798 53648 239120 53928
rect 798 53248 239200 53648
rect 798 52968 239120 53248
rect 798 52568 239200 52968
rect 798 52288 239120 52568
rect 798 51888 239200 52288
rect 798 51608 239120 51888
rect 798 51208 239200 51608
rect 798 50928 239120 51208
rect 798 50528 239200 50928
rect 798 50248 239120 50528
rect 798 49848 239200 50248
rect 798 49568 239120 49848
rect 798 49168 239200 49568
rect 798 48888 239120 49168
rect 798 48488 239200 48888
rect 798 48208 239120 48488
rect 798 47808 239200 48208
rect 798 47528 239120 47808
rect 798 47128 239200 47528
rect 798 46848 239120 47128
rect 798 46448 239200 46848
rect 798 46168 239120 46448
rect 798 45768 239200 46168
rect 798 45488 239120 45768
rect 798 2143 239200 45488
<< metal4 >>
rect -1076 -4 -756 199652
rect -416 656 -96 198992
rect 4208 -4 4528 199652
rect 4868 -4 5188 199652
rect 34928 172874 35248 199652
rect 35588 172874 35908 199652
rect 65648 172874 65968 199652
rect 66308 172874 66628 199652
rect 34928 72874 35248 119864
rect 35588 72874 35908 119680
rect 65648 72874 65968 119864
rect 66308 72874 66628 119864
rect 34928 -4 35248 19864
rect 35588 -4 35908 19680
rect 65648 -4 65968 19864
rect 66308 -4 66628 19864
rect 96368 -4 96688 199652
rect 97028 -4 97348 199652
rect 127088 -4 127408 199652
rect 127748 -4 128068 199652
rect 157808 172874 158128 199652
rect 158468 172874 158788 199652
rect 188528 172874 188848 199652
rect 189188 172874 189508 199652
rect 157808 72874 158128 119680
rect 158468 72874 158788 119864
rect 188528 72874 188848 119864
rect 189188 72874 189508 119864
rect 157808 -4 158128 19680
rect 158468 -4 158788 19864
rect 188528 -4 188848 19864
rect 189188 -4 189508 19864
rect 219248 -4 219568 199652
rect 219908 -4 220228 199652
rect 240032 656 240352 198992
rect 240692 -4 241012 199652
<< obsm4 >>
rect 17723 172794 34848 197165
rect 35328 172794 35508 197165
rect 35988 172794 65568 197165
rect 66048 172794 66228 197165
rect 66708 172794 96288 197165
rect 17723 119944 96288 172794
rect 17723 72794 34848 119944
rect 35328 119760 65568 119944
rect 35328 72794 35508 119760
rect 35988 72794 65568 119760
rect 66048 72794 66228 119944
rect 66708 72794 96288 119944
rect 17723 19944 96288 72794
rect 17723 17035 34848 19944
rect 35328 19760 65568 19944
rect 35328 17035 35508 19760
rect 35988 17035 65568 19760
rect 66048 17035 66228 19944
rect 66708 17035 96288 19944
rect 96768 17035 96948 197165
rect 97428 17035 127008 197165
rect 127488 17035 127668 197165
rect 128148 172794 157728 197165
rect 158208 172794 158388 197165
rect 158868 172794 188448 197165
rect 188928 172794 189108 197165
rect 189588 172794 209149 197165
rect 128148 119944 209149 172794
rect 128148 119760 158388 119944
rect 128148 72794 157728 119760
rect 158208 72794 158388 119760
rect 158868 72794 188448 119944
rect 188928 72794 189108 119944
rect 189588 72794 209149 119944
rect 128148 19944 209149 72794
rect 128148 19760 158388 19944
rect 128148 17035 157728 19760
rect 158208 17035 158388 19760
rect 158868 17035 188448 19944
rect 188928 17035 189108 19944
rect 189588 17035 209149 19944
<< metal5 >>
rect -1076 199332 241012 199652
rect -416 198672 240352 198992
rect -1076 189822 241012 190142
rect -1076 189162 241012 189482
rect -1076 159186 241012 159506
rect -1076 158526 241012 158846
rect -1076 128550 241012 128870
rect -1076 127890 241012 128210
rect -1076 97914 241012 98234
rect -1076 97254 241012 97574
rect -1076 67278 241012 67598
rect -1076 66618 241012 66938
rect -1076 36642 241012 36962
rect -1076 35982 241012 36302
rect -1076 6006 241012 6326
rect -1076 5346 241012 5666
rect -416 656 240352 976
rect -1076 -4 241012 316
<< obsm5 >>
rect 19068 159826 160516 174580
rect 19068 129190 160516 158206
rect 19068 98554 160516 127570
rect 19068 67918 160516 96934
rect 19068 37282 160516 66298
rect 19068 17180 160516 35662
<< labels >>
rlabel metal2 s 26422 0 26478 800 6 clk
port 1 nsew signal input
rlabel metal3 s 239200 45568 240000 45688 6 in_data[0]
port 2 nsew signal input
rlabel metal3 s 239200 110168 240000 110288 6 in_data[100]
port 3 nsew signal input
rlabel metal3 s 239200 53048 240000 53168 6 in_data[101]
port 4 nsew signal input
rlabel metal3 s 239200 53728 240000 53848 6 in_data[102]
port 5 nsew signal input
rlabel metal3 s 239200 55088 240000 55208 6 in_data[103]
port 6 nsew signal input
rlabel metal3 s 239200 57128 240000 57248 6 in_data[104]
port 7 nsew signal input
rlabel metal3 s 239200 58488 240000 58608 6 in_data[105]
port 8 nsew signal input
rlabel metal3 s 239200 56448 240000 56568 6 in_data[106]
port 9 nsew signal input
rlabel metal3 s 239200 109488 240000 109608 6 in_data[107]
port 10 nsew signal input
rlabel metal3 s 239200 108128 240000 108248 6 in_data[108]
port 11 nsew signal input
rlabel metal3 s 239200 87728 240000 87848 6 in_data[109]
port 12 nsew signal input
rlabel metal3 s 239200 61208 240000 61328 6 in_data[10]
port 13 nsew signal input
rlabel metal3 s 239200 101328 240000 101448 6 in_data[110]
port 14 nsew signal input
rlabel metal3 s 239200 52368 240000 52488 6 in_data[111]
port 15 nsew signal input
rlabel metal3 s 239200 106088 240000 106208 6 in_data[112]
port 16 nsew signal input
rlabel metal3 s 239200 104728 240000 104848 6 in_data[113]
port 17 nsew signal input
rlabel metal3 s 239200 105408 240000 105528 6 in_data[114]
port 18 nsew signal input
rlabel metal3 s 239200 107448 240000 107568 6 in_data[115]
port 19 nsew signal input
rlabel metal3 s 239200 99288 240000 99408 6 in_data[116]
port 20 nsew signal input
rlabel metal2 s 149426 199200 149482 200000 6 in_data[117]
port 21 nsew signal input
rlabel metal2 s 141054 199200 141110 200000 6 in_data[118]
port 22 nsew signal input
rlabel metal2 s 144918 199200 144974 200000 6 in_data[119]
port 23 nsew signal input
rlabel metal3 s 239200 46248 240000 46368 6 in_data[11]
port 24 nsew signal input
rlabel metal2 s 155222 199200 155278 200000 6 in_data[120]
port 25 nsew signal input
rlabel metal2 s 150714 199200 150770 200000 6 in_data[121]
port 26 nsew signal input
rlabel metal2 s 154578 199200 154634 200000 6 in_data[122]
port 27 nsew signal input
rlabel metal2 s 168102 199200 168158 200000 6 in_data[123]
port 28 nsew signal input
rlabel metal2 s 164882 199200 164938 200000 6 in_data[124]
port 29 nsew signal input
rlabel metal2 s 163594 199200 163650 200000 6 in_data[125]
port 30 nsew signal input
rlabel metal2 s 152002 199200 152058 200000 6 in_data[126]
port 31 nsew signal input
rlabel metal3 s 239200 89088 240000 89208 6 in_data[127]
port 32 nsew signal input
rlabel metal3 s 239200 85688 240000 85808 6 in_data[12]
port 33 nsew signal input
rlabel metal3 s 239200 83648 240000 83768 6 in_data[13]
port 34 nsew signal input
rlabel metal3 s 239200 87048 240000 87168 6 in_data[14]
port 35 nsew signal input
rlabel metal3 s 239200 82968 240000 83088 6 in_data[15]
port 36 nsew signal input
rlabel metal3 s 239200 98608 240000 98728 6 in_data[16]
port 37 nsew signal input
rlabel metal3 s 239200 96568 240000 96688 6 in_data[17]
port 38 nsew signal input
rlabel metal3 s 239200 97928 240000 98048 6 in_data[18]
port 39 nsew signal input
rlabel metal3 s 239200 99968 240000 100088 6 in_data[19]
port 40 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 in_data[1]
port 41 nsew signal input
rlabel metal3 s 239200 106768 240000 106888 6 in_data[20]
port 42 nsew signal input
rlabel metal2 s 135258 199200 135314 200000 6 in_data[21]
port 43 nsew signal input
rlabel metal2 s 146850 199200 146906 200000 6 in_data[22]
port 44 nsew signal input
rlabel metal2 s 138478 199200 138534 200000 6 in_data[23]
port 45 nsew signal input
rlabel metal2 s 160374 199200 160430 200000 6 in_data[24]
port 46 nsew signal input
rlabel metal2 s 161018 199200 161074 200000 6 in_data[25]
port 47 nsew signal input
rlabel metal2 s 159730 199200 159786 200000 6 in_data[26]
port 48 nsew signal input
rlabel metal2 s 162950 199200 163006 200000 6 in_data[27]
port 49 nsew signal input
rlabel metal2 s 161662 199200 161718 200000 6 in_data[28]
port 50 nsew signal input
rlabel metal2 s 162306 199200 162362 200000 6 in_data[29]
port 51 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 in_data[2]
port 52 nsew signal input
rlabel metal2 s 159086 199200 159142 200000 6 in_data[30]
port 53 nsew signal input
rlabel metal2 s 148138 199200 148194 200000 6 in_data[31]
port 54 nsew signal input
rlabel metal3 s 239200 70048 240000 70168 6 in_data[32]
port 55 nsew signal input
rlabel metal3 s 239200 59848 240000 59968 6 in_data[33]
port 56 nsew signal input
rlabel metal3 s 239200 63248 240000 63368 6 in_data[34]
port 57 nsew signal input
rlabel metal3 s 239200 64608 240000 64728 6 in_data[35]
port 58 nsew signal input
rlabel metal3 s 239200 78208 240000 78328 6 in_data[36]
port 59 nsew signal input
rlabel metal3 s 239200 54408 240000 54528 6 in_data[37]
port 60 nsew signal input
rlabel metal3 s 239200 68688 240000 68808 6 in_data[38]
port 61 nsew signal input
rlabel metal3 s 239200 70728 240000 70848 6 in_data[39]
port 62 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 in_data[3]
port 63 nsew signal input
rlabel metal3 s 239200 61888 240000 62008 6 in_data[40]
port 64 nsew signal input
rlabel metal3 s 239200 66648 240000 66768 6 in_data[41]
port 65 nsew signal input
rlabel metal3 s 239200 72768 240000 72888 6 in_data[42]
port 66 nsew signal input
rlabel metal3 s 239200 82288 240000 82408 6 in_data[43]
port 67 nsew signal input
rlabel metal3 s 239200 79568 240000 79688 6 in_data[44]
port 68 nsew signal input
rlabel metal3 s 239200 85008 240000 85128 6 in_data[45]
port 69 nsew signal input
rlabel metal3 s 239200 94528 240000 94648 6 in_data[46]
port 70 nsew signal input
rlabel metal3 s 239200 74808 240000 74928 6 in_data[47]
port 71 nsew signal input
rlabel metal3 s 239200 93848 240000 93968 6 in_data[48]
port 72 nsew signal input
rlabel metal3 s 239200 91808 240000 91928 6 in_data[49]
port 73 nsew signal input
rlabel metal3 s 239200 67328 240000 67448 6 in_data[4]
port 74 nsew signal input
rlabel metal3 s 239200 91128 240000 91248 6 in_data[50]
port 75 nsew signal input
rlabel metal3 s 239200 93168 240000 93288 6 in_data[51]
port 76 nsew signal input
rlabel metal3 s 239200 95208 240000 95328 6 in_data[52]
port 77 nsew signal input
rlabel metal2 s 139766 199200 139822 200000 6 in_data[53]
port 78 nsew signal input
rlabel metal2 s 143630 199200 143686 200000 6 in_data[54]
port 79 nsew signal input
rlabel metal2 s 144274 199200 144330 200000 6 in_data[55]
port 80 nsew signal input
rlabel metal2 s 165526 199200 165582 200000 6 in_data[56]
port 81 nsew signal input
rlabel metal2 s 166170 199200 166226 200000 6 in_data[57]
port 82 nsew signal input
rlabel metal2 s 166814 199200 166870 200000 6 in_data[58]
port 83 nsew signal input
rlabel metal2 s 157154 199200 157210 200000 6 in_data[59]
port 84 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 in_data[5]
port 85 nsew signal input
rlabel metal2 s 158442 199200 158498 200000 6 in_data[60]
port 86 nsew signal input
rlabel metal2 s 157798 199200 157854 200000 6 in_data[61]
port 87 nsew signal input
rlabel metal2 s 155866 199200 155922 200000 6 in_data[62]
port 88 nsew signal input
rlabel metal3 s 239200 102688 240000 102808 6 in_data[63]
port 89 nsew signal input
rlabel metal3 s 239200 72088 240000 72208 6 in_data[64]
port 90 nsew signal input
rlabel metal3 s 239200 59168 240000 59288 6 in_data[65]
port 91 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 in_data[66]
port 92 nsew signal input
rlabel metal3 s 239200 60528 240000 60648 6 in_data[67]
port 93 nsew signal input
rlabel metal3 s 239200 73448 240000 73568 6 in_data[68]
port 94 nsew signal input
rlabel metal3 s 239200 65288 240000 65408 6 in_data[69]
port 95 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 in_data[6]
port 96 nsew signal input
rlabel metal3 s 239200 68008 240000 68128 6 in_data[70]
port 97 nsew signal input
rlabel metal3 s 239200 69368 240000 69488 6 in_data[71]
port 98 nsew signal input
rlabel metal3 s 239200 62568 240000 62688 6 in_data[72]
port 99 nsew signal input
rlabel metal3 s 239200 57808 240000 57928 6 in_data[73]
port 100 nsew signal input
rlabel metal3 s 239200 55768 240000 55888 6 in_data[74]
port 101 nsew signal input
rlabel metal3 s 239200 84328 240000 84448 6 in_data[75]
port 102 nsew signal input
rlabel metal3 s 239200 78888 240000 79008 6 in_data[76]
port 103 nsew signal input
rlabel metal3 s 239200 86368 240000 86488 6 in_data[77]
port 104 nsew signal input
rlabel metal3 s 239200 88408 240000 88528 6 in_data[78]
port 105 nsew signal input
rlabel metal3 s 239200 47608 240000 47728 6 in_data[79]
port 106 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 in_data[7]
port 107 nsew signal input
rlabel metal3 s 239200 95888 240000 96008 6 in_data[80]
port 108 nsew signal input
rlabel metal3 s 239200 100648 240000 100768 6 in_data[81]
port 109 nsew signal input
rlabel metal3 s 239200 92488 240000 92608 6 in_data[82]
port 110 nsew signal input
rlabel metal3 s 239200 104048 240000 104168 6 in_data[83]
port 111 nsew signal input
rlabel metal3 s 239200 97248 240000 97368 6 in_data[84]
port 112 nsew signal input
rlabel metal2 s 139122 199200 139178 200000 6 in_data[85]
port 113 nsew signal input
rlabel metal2 s 140410 199200 140466 200000 6 in_data[86]
port 114 nsew signal input
rlabel metal2 s 142986 199200 143042 200000 6 in_data[87]
port 115 nsew signal input
rlabel metal2 s 151358 199200 151414 200000 6 in_data[88]
port 116 nsew signal input
rlabel metal2 s 152646 199200 152702 200000 6 in_data[89]
port 117 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 in_data[8]
port 118 nsew signal input
rlabel metal2 s 153934 199200 153990 200000 6 in_data[90]
port 119 nsew signal input
rlabel metal2 s 167458 199200 167514 200000 6 in_data[91]
port 120 nsew signal input
rlabel metal2 s 156510 199200 156566 200000 6 in_data[92]
port 121 nsew signal input
rlabel metal2 s 164238 199200 164294 200000 6 in_data[93]
port 122 nsew signal input
rlabel metal2 s 153290 199200 153346 200000 6 in_data[94]
port 123 nsew signal input
rlabel metal3 s 239200 89768 240000 89888 6 in_data[95]
port 124 nsew signal input
rlabel metal3 s 239200 71408 240000 71528 6 in_data[96]
port 125 nsew signal input
rlabel metal3 s 239200 65968 240000 66088 6 in_data[97]
port 126 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 in_data[98]
port 127 nsew signal input
rlabel metal3 s 239200 63928 240000 64048 6 in_data[99]
port 128 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 in_data[9]
port 129 nsew signal input
rlabel metal3 s 239200 103368 240000 103488 6 in_ready
port 130 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 out_data[0]
port 131 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 out_data[100]
port 132 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 out_data[101]
port 133 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 out_data[102]
port 134 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 out_data[103]
port 135 nsew signal output
rlabel metal3 s 239200 80248 240000 80368 6 out_data[104]
port 136 nsew signal output
rlabel metal3 s 239200 46928 240000 47048 6 out_data[105]
port 137 nsew signal output
rlabel metal3 s 239200 51008 240000 51128 6 out_data[106]
port 138 nsew signal output
rlabel metal3 s 239200 48288 240000 48408 6 out_data[107]
port 139 nsew signal output
rlabel metal3 s 239200 90448 240000 90568 6 out_data[108]
port 140 nsew signal output
rlabel metal2 s 112718 199200 112774 200000 6 out_data[109]
port 141 nsew signal output
rlabel metal3 s 239200 50328 240000 50448 6 out_data[10]
port 142 nsew signal output
rlabel metal2 s 117870 199200 117926 200000 6 out_data[110]
port 143 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 out_data[111]
port 144 nsew signal output
rlabel metal2 s 95330 199200 95386 200000 6 out_data[112]
port 145 nsew signal output
rlabel metal2 s 93398 199200 93454 200000 6 out_data[113]
port 146 nsew signal output
rlabel metal2 s 92754 199200 92810 200000 6 out_data[114]
port 147 nsew signal output
rlabel metal2 s 87602 199200 87658 200000 6 out_data[115]
port 148 nsew signal output
rlabel metal2 s 89534 199200 89590 200000 6 out_data[116]
port 149 nsew signal output
rlabel metal2 s 90822 199200 90878 200000 6 out_data[117]
port 150 nsew signal output
rlabel metal2 s 92110 199200 92166 200000 6 out_data[118]
port 151 nsew signal output
rlabel metal2 s 104990 199200 105046 200000 6 out_data[119]
port 152 nsew signal output
rlabel metal3 s 239200 76848 240000 76968 6 out_data[11]
port 153 nsew signal output
rlabel metal2 s 137834 199200 137890 200000 6 out_data[120]
port 154 nsew signal output
rlabel metal2 s 145562 199200 145618 200000 6 out_data[121]
port 155 nsew signal output
rlabel metal2 s 137190 199200 137246 200000 6 out_data[122]
port 156 nsew signal output
rlabel metal2 s 147494 199200 147550 200000 6 out_data[123]
port 157 nsew signal output
rlabel metal2 s 134614 199200 134670 200000 6 out_data[124]
port 158 nsew signal output
rlabel metal2 s 135902 199200 135958 200000 6 out_data[125]
port 159 nsew signal output
rlabel metal2 s 129462 199200 129518 200000 6 out_data[126]
port 160 nsew signal output
rlabel metal2 s 124310 199200 124366 200000 6 out_data[127]
port 161 nsew signal output
rlabel metal2 s 117226 199200 117282 200000 6 out_data[12]
port 162 nsew signal output
rlabel metal2 s 123666 199200 123722 200000 6 out_data[13]
port 163 nsew signal output
rlabel metal2 s 124954 199200 125010 200000 6 out_data[14]
port 164 nsew signal output
rlabel metal2 s 119158 199200 119214 200000 6 out_data[15]
port 165 nsew signal output
rlabel metal2 s 102414 199200 102470 200000 6 out_data[16]
port 166 nsew signal output
rlabel metal2 s 97262 199200 97318 200000 6 out_data[17]
port 167 nsew signal output
rlabel metal2 s 94686 199200 94742 200000 6 out_data[18]
port 168 nsew signal output
rlabel metal2 s 94042 199200 94098 200000 6 out_data[19]
port 169 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 out_data[1]
port 170 nsew signal output
rlabel metal2 s 91466 199200 91522 200000 6 out_data[20]
port 171 nsew signal output
rlabel metal2 s 90178 199200 90234 200000 6 out_data[21]
port 172 nsew signal output
rlabel metal2 s 101770 199200 101826 200000 6 out_data[22]
port 173 nsew signal output
rlabel metal2 s 104346 199200 104402 200000 6 out_data[23]
port 174 nsew signal output
rlabel metal2 s 146206 199200 146262 200000 6 out_data[24]
port 175 nsew signal output
rlabel metal2 s 148782 199200 148838 200000 6 out_data[25]
port 176 nsew signal output
rlabel metal2 s 115938 199200 115994 200000 6 out_data[26]
port 177 nsew signal output
rlabel metal2 s 133326 199200 133382 200000 6 out_data[27]
port 178 nsew signal output
rlabel metal2 s 114006 199200 114062 200000 6 out_data[28]
port 179 nsew signal output
rlabel metal2 s 126242 199200 126298 200000 6 out_data[29]
port 180 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 out_data[2]
port 181 nsew signal output
rlabel metal2 s 123022 199200 123078 200000 6 out_data[30]
port 182 nsew signal output
rlabel metal2 s 114650 199200 114706 200000 6 out_data[31]
port 183 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 out_data[32]
port 184 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 out_data[33]
port 185 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 out_data[34]
port 186 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 out_data[35]
port 187 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 out_data[36]
port 188 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 out_data[37]
port 189 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 out_data[38]
port 190 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 out_data[39]
port 191 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 out_data[3]
port 192 nsew signal output
rlabel metal3 s 239200 81608 240000 81728 6 out_data[40]
port 193 nsew signal output
rlabel metal3 s 239200 76168 240000 76288 6 out_data[41]
port 194 nsew signal output
rlabel metal3 s 239200 51688 240000 51808 6 out_data[42]
port 195 nsew signal output
rlabel metal3 s 239200 49648 240000 49768 6 out_data[43]
port 196 nsew signal output
rlabel metal2 s 113362 199200 113418 200000 6 out_data[44]
port 197 nsew signal output
rlabel metal2 s 127530 199200 127586 200000 6 out_data[45]
port 198 nsew signal output
rlabel metal2 s 120446 199200 120502 200000 6 out_data[46]
port 199 nsew signal output
rlabel metal2 s 121734 199200 121790 200000 6 out_data[47]
port 200 nsew signal output
rlabel metal2 s 98550 199200 98606 200000 6 out_data[48]
port 201 nsew signal output
rlabel metal2 s 99194 199200 99250 200000 6 out_data[49]
port 202 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 out_data[4]
port 203 nsew signal output
rlabel metal2 s 99838 199200 99894 200000 6 out_data[50]
port 204 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 out_data[51]
port 205 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 out_data[52]
port 206 nsew signal output
rlabel metal2 s 88890 199200 88946 200000 6 out_data[53]
port 207 nsew signal output
rlabel metal2 s 100482 199200 100538 200000 6 out_data[54]
port 208 nsew signal output
rlabel metal2 s 103702 199200 103758 200000 6 out_data[55]
port 209 nsew signal output
rlabel metal2 s 141698 199200 141754 200000 6 out_data[56]
port 210 nsew signal output
rlabel metal2 s 132682 199200 132738 200000 6 out_data[57]
port 211 nsew signal output
rlabel metal2 s 125598 199200 125654 200000 6 out_data[58]
port 212 nsew signal output
rlabel metal2 s 133970 199200 134026 200000 6 out_data[59]
port 213 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 out_data[5]
port 214 nsew signal output
rlabel metal2 s 128818 199200 128874 200000 6 out_data[60]
port 215 nsew signal output
rlabel metal2 s 116582 199200 116638 200000 6 out_data[61]
port 216 nsew signal output
rlabel metal2 s 130106 199200 130162 200000 6 out_data[62]
port 217 nsew signal output
rlabel metal2 s 115294 199200 115350 200000 6 out_data[63]
port 218 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 out_data[64]
port 219 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 out_data[65]
port 220 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 out_data[66]
port 221 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 out_data[67]
port 222 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 out_data[68]
port 223 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 out_data[69]
port 224 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 out_data[6]
port 225 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 out_data[70]
port 226 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 out_data[71]
port 227 nsew signal output
rlabel metal3 s 239200 80928 240000 81048 6 out_data[72]
port 228 nsew signal output
rlabel metal3 s 239200 75488 240000 75608 6 out_data[73]
port 229 nsew signal output
rlabel metal3 s 239200 74128 240000 74248 6 out_data[74]
port 230 nsew signal output
rlabel metal3 s 239200 48968 240000 49088 6 out_data[75]
port 231 nsew signal output
rlabel metal2 s 126886 199200 126942 200000 6 out_data[76]
port 232 nsew signal output
rlabel metal2 s 121090 199200 121146 200000 6 out_data[77]
port 233 nsew signal output
rlabel metal2 s 118514 199200 118570 200000 6 out_data[78]
port 234 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 out_data[79]
port 235 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 out_data[7]
port 236 nsew signal output
rlabel metal2 s 97906 199200 97962 200000 6 out_data[80]
port 237 nsew signal output
rlabel metal2 s 95974 199200 96030 200000 6 out_data[81]
port 238 nsew signal output
rlabel metal2 s 96618 199200 96674 200000 6 out_data[82]
port 239 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 out_data[83]
port 240 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 out_data[84]
port 241 nsew signal output
rlabel metal2 s 88246 199200 88302 200000 6 out_data[85]
port 242 nsew signal output
rlabel metal2 s 101126 199200 101182 200000 6 out_data[86]
port 243 nsew signal output
rlabel metal2 s 103058 199200 103114 200000 6 out_data[87]
port 244 nsew signal output
rlabel metal2 s 142342 199200 142398 200000 6 out_data[88]
port 245 nsew signal output
rlabel metal2 s 131394 199200 131450 200000 6 out_data[89]
port 246 nsew signal output
rlabel metal3 s 239200 108808 240000 108928 6 out_data[8]
port 247 nsew signal output
rlabel metal2 s 150070 199200 150126 200000 6 out_data[90]
port 248 nsew signal output
rlabel metal2 s 136546 199200 136602 200000 6 out_data[91]
port 249 nsew signal output
rlabel metal2 s 130750 199200 130806 200000 6 out_data[92]
port 250 nsew signal output
rlabel metal2 s 132038 199200 132094 200000 6 out_data[93]
port 251 nsew signal output
rlabel metal2 s 128174 199200 128230 200000 6 out_data[94]
port 252 nsew signal output
rlabel metal2 s 119802 199200 119858 200000 6 out_data[95]
port 253 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 out_data[96]
port 254 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 out_data[97]
port 255 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 out_data[98]
port 256 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 out_data[99]
port 257 nsew signal output
rlabel metal3 s 239200 77528 240000 77648 6 out_data[9]
port 258 nsew signal output
rlabel metal2 s 122378 199200 122434 200000 6 out_ready
port 259 nsew signal output
rlabel metal3 s 239200 102008 240000 102128 6 reset
port 260 nsew signal input
rlabel metal2 s 207386 199200 207442 200000 6 s_box_ready
port 261 nsew signal output
rlabel metal4 s -416 656 -96 198992 4 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -416 656 240352 976 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -416 198672 240352 198992 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 240032 656 240352 198992 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 4208 -4 4528 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 34928 -4 35248 19864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 34928 72874 35248 119864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 34928 172874 35248 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 65648 -4 65968 19864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 65648 72874 65968 119864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 65648 172874 65968 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 96368 -4 96688 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 127088 -4 127408 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 157808 -4 158128 19680 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 157808 72874 158128 119680 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 157808 172874 158128 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 188528 -4 188848 19864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 188528 72874 188848 119864 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 188528 172874 188848 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s 219248 -4 219568 199652 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 5346 241012 5666 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 35982 241012 36302 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 66618 241012 66938 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 97254 241012 97574 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 127890 241012 128210 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 158526 241012 158846 6 vccd1
port 262 nsew power bidirectional
rlabel metal5 s -1076 189162 241012 189482 6 vccd1
port 262 nsew power bidirectional
rlabel metal4 s -1076 -4 -756 199652 4 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 -4 241012 316 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 199332 241012 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 240692 -4 241012 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 4868 -4 5188 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 35588 -4 35908 19680 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 35588 72874 35908 119680 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 35588 172874 35908 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 66308 -4 66628 19864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 66308 72874 66628 119864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 66308 172874 66628 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 97028 -4 97348 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 127748 -4 128068 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 158468 -4 158788 19864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 158468 72874 158788 119864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 158468 172874 158788 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 189188 -4 189508 19864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 189188 72874 189508 119864 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 189188 172874 189508 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal4 s 219908 -4 220228 199652 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 6006 241012 6326 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 36642 241012 36962 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 67278 241012 67598 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 97914 241012 98234 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 128550 241012 128870 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 159186 241012 159506 6 vssd1
port 263 nsew ground bidirectional
rlabel metal5 s -1076 189822 241012 190142 6 vssd1
port 263 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 240000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16931310
string GDS_FILE /openlane/designs/subBytes_asic/runs/full_guide/results/signoff/subBytes_asic.magic.gds
string GDS_START 6569284
<< end >>

