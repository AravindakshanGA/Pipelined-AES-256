magic
tech sky130A
magscale 1 2
timestamp 1543373562
<< checkpaint >>
rect -1302 -1365 21270 26645
<< metal1 >>
rect 78 0 114 25280
rect 150 0 186 25280
rect 222 24569 258 25201
rect 222 23779 258 24411
rect 222 22989 258 23621
rect 222 22199 258 22831
rect 222 21409 258 22041
rect 222 20619 258 21251
rect 222 19829 258 20461
rect 222 19039 258 19671
rect 222 18249 258 18881
rect 222 17459 258 18091
rect 222 16669 258 17301
rect 222 15879 258 16511
rect 222 15089 258 15721
rect 222 14299 258 14931
rect 222 13509 258 14141
rect 222 12719 258 13351
rect 222 11929 258 12561
rect 222 11139 258 11771
rect 222 10349 258 10981
rect 222 9559 258 10191
rect 222 8769 258 9401
rect 222 7979 258 8611
rect 222 7189 258 7821
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 79 258 711
rect 294 0 330 25280
rect 366 0 402 25280
rect 846 0 882 25280
rect 918 0 954 25280
rect 990 24569 1026 25201
rect 990 23779 1026 24411
rect 990 22989 1026 23621
rect 990 22199 1026 22831
rect 990 21409 1026 22041
rect 990 20619 1026 21251
rect 990 19829 1026 20461
rect 990 19039 1026 19671
rect 990 18249 1026 18881
rect 990 17459 1026 18091
rect 990 16669 1026 17301
rect 990 15879 1026 16511
rect 990 15089 1026 15721
rect 990 14299 1026 14931
rect 990 13509 1026 14141
rect 990 12719 1026 13351
rect 990 11929 1026 12561
rect 990 11139 1026 11771
rect 990 10349 1026 10981
rect 990 9559 1026 10191
rect 990 8769 1026 9401
rect 990 7979 1026 8611
rect 990 7189 1026 7821
rect 990 6399 1026 7031
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 79 1026 711
rect 1062 0 1098 25280
rect 1134 0 1170 25280
rect 1326 0 1362 25280
rect 1398 0 1434 25280
rect 1470 24569 1506 25201
rect 1470 23779 1506 24411
rect 1470 22989 1506 23621
rect 1470 22199 1506 22831
rect 1470 21409 1506 22041
rect 1470 20619 1506 21251
rect 1470 19829 1506 20461
rect 1470 19039 1506 19671
rect 1470 18249 1506 18881
rect 1470 17459 1506 18091
rect 1470 16669 1506 17301
rect 1470 15879 1506 16511
rect 1470 15089 1506 15721
rect 1470 14299 1506 14931
rect 1470 13509 1506 14141
rect 1470 12719 1506 13351
rect 1470 11929 1506 12561
rect 1470 11139 1506 11771
rect 1470 10349 1506 10981
rect 1470 9559 1506 10191
rect 1470 8769 1506 9401
rect 1470 7979 1506 8611
rect 1470 7189 1506 7821
rect 1470 6399 1506 7031
rect 1470 5609 1506 6241
rect 1470 4819 1506 5451
rect 1470 4029 1506 4661
rect 1470 3239 1506 3871
rect 1470 2449 1506 3081
rect 1470 1659 1506 2291
rect 1470 869 1506 1501
rect 1470 79 1506 711
rect 1542 0 1578 25280
rect 1614 0 1650 25280
rect 2094 0 2130 25280
rect 2166 0 2202 25280
rect 2238 24569 2274 25201
rect 2238 23779 2274 24411
rect 2238 22989 2274 23621
rect 2238 22199 2274 22831
rect 2238 21409 2274 22041
rect 2238 20619 2274 21251
rect 2238 19829 2274 20461
rect 2238 19039 2274 19671
rect 2238 18249 2274 18881
rect 2238 17459 2274 18091
rect 2238 16669 2274 17301
rect 2238 15879 2274 16511
rect 2238 15089 2274 15721
rect 2238 14299 2274 14931
rect 2238 13509 2274 14141
rect 2238 12719 2274 13351
rect 2238 11929 2274 12561
rect 2238 11139 2274 11771
rect 2238 10349 2274 10981
rect 2238 9559 2274 10191
rect 2238 8769 2274 9401
rect 2238 7979 2274 8611
rect 2238 7189 2274 7821
rect 2238 6399 2274 7031
rect 2238 5609 2274 6241
rect 2238 4819 2274 5451
rect 2238 4029 2274 4661
rect 2238 3239 2274 3871
rect 2238 2449 2274 3081
rect 2238 1659 2274 2291
rect 2238 869 2274 1501
rect 2238 79 2274 711
rect 2310 0 2346 25280
rect 2382 0 2418 25280
rect 2574 0 2610 25280
rect 2646 0 2682 25280
rect 2718 24569 2754 25201
rect 2718 23779 2754 24411
rect 2718 22989 2754 23621
rect 2718 22199 2754 22831
rect 2718 21409 2754 22041
rect 2718 20619 2754 21251
rect 2718 19829 2754 20461
rect 2718 19039 2754 19671
rect 2718 18249 2754 18881
rect 2718 17459 2754 18091
rect 2718 16669 2754 17301
rect 2718 15879 2754 16511
rect 2718 15089 2754 15721
rect 2718 14299 2754 14931
rect 2718 13509 2754 14141
rect 2718 12719 2754 13351
rect 2718 11929 2754 12561
rect 2718 11139 2754 11771
rect 2718 10349 2754 10981
rect 2718 9559 2754 10191
rect 2718 8769 2754 9401
rect 2718 7979 2754 8611
rect 2718 7189 2754 7821
rect 2718 6399 2754 7031
rect 2718 5609 2754 6241
rect 2718 4819 2754 5451
rect 2718 4029 2754 4661
rect 2718 3239 2754 3871
rect 2718 2449 2754 3081
rect 2718 1659 2754 2291
rect 2718 869 2754 1501
rect 2718 79 2754 711
rect 2790 0 2826 25280
rect 2862 0 2898 25280
rect 3342 0 3378 25280
rect 3414 0 3450 25280
rect 3486 24569 3522 25201
rect 3486 23779 3522 24411
rect 3486 22989 3522 23621
rect 3486 22199 3522 22831
rect 3486 21409 3522 22041
rect 3486 20619 3522 21251
rect 3486 19829 3522 20461
rect 3486 19039 3522 19671
rect 3486 18249 3522 18881
rect 3486 17459 3522 18091
rect 3486 16669 3522 17301
rect 3486 15879 3522 16511
rect 3486 15089 3522 15721
rect 3486 14299 3522 14931
rect 3486 13509 3522 14141
rect 3486 12719 3522 13351
rect 3486 11929 3522 12561
rect 3486 11139 3522 11771
rect 3486 10349 3522 10981
rect 3486 9559 3522 10191
rect 3486 8769 3522 9401
rect 3486 7979 3522 8611
rect 3486 7189 3522 7821
rect 3486 6399 3522 7031
rect 3486 5609 3522 6241
rect 3486 4819 3522 5451
rect 3486 4029 3522 4661
rect 3486 3239 3522 3871
rect 3486 2449 3522 3081
rect 3486 1659 3522 2291
rect 3486 869 3522 1501
rect 3486 79 3522 711
rect 3558 0 3594 25280
rect 3630 0 3666 25280
rect 3822 0 3858 25280
rect 3894 0 3930 25280
rect 3966 24569 4002 25201
rect 3966 23779 4002 24411
rect 3966 22989 4002 23621
rect 3966 22199 4002 22831
rect 3966 21409 4002 22041
rect 3966 20619 4002 21251
rect 3966 19829 4002 20461
rect 3966 19039 4002 19671
rect 3966 18249 4002 18881
rect 3966 17459 4002 18091
rect 3966 16669 4002 17301
rect 3966 15879 4002 16511
rect 3966 15089 4002 15721
rect 3966 14299 4002 14931
rect 3966 13509 4002 14141
rect 3966 12719 4002 13351
rect 3966 11929 4002 12561
rect 3966 11139 4002 11771
rect 3966 10349 4002 10981
rect 3966 9559 4002 10191
rect 3966 8769 4002 9401
rect 3966 7979 4002 8611
rect 3966 7189 4002 7821
rect 3966 6399 4002 7031
rect 3966 5609 4002 6241
rect 3966 4819 4002 5451
rect 3966 4029 4002 4661
rect 3966 3239 4002 3871
rect 3966 2449 4002 3081
rect 3966 1659 4002 2291
rect 3966 869 4002 1501
rect 3966 79 4002 711
rect 4038 0 4074 25280
rect 4110 0 4146 25280
rect 4590 0 4626 25280
rect 4662 0 4698 25280
rect 4734 24569 4770 25201
rect 4734 23779 4770 24411
rect 4734 22989 4770 23621
rect 4734 22199 4770 22831
rect 4734 21409 4770 22041
rect 4734 20619 4770 21251
rect 4734 19829 4770 20461
rect 4734 19039 4770 19671
rect 4734 18249 4770 18881
rect 4734 17459 4770 18091
rect 4734 16669 4770 17301
rect 4734 15879 4770 16511
rect 4734 15089 4770 15721
rect 4734 14299 4770 14931
rect 4734 13509 4770 14141
rect 4734 12719 4770 13351
rect 4734 11929 4770 12561
rect 4734 11139 4770 11771
rect 4734 10349 4770 10981
rect 4734 9559 4770 10191
rect 4734 8769 4770 9401
rect 4734 7979 4770 8611
rect 4734 7189 4770 7821
rect 4734 6399 4770 7031
rect 4734 5609 4770 6241
rect 4734 4819 4770 5451
rect 4734 4029 4770 4661
rect 4734 3239 4770 3871
rect 4734 2449 4770 3081
rect 4734 1659 4770 2291
rect 4734 869 4770 1501
rect 4734 79 4770 711
rect 4806 0 4842 25280
rect 4878 0 4914 25280
rect 5070 0 5106 25280
rect 5142 0 5178 25280
rect 5214 24569 5250 25201
rect 5214 23779 5250 24411
rect 5214 22989 5250 23621
rect 5214 22199 5250 22831
rect 5214 21409 5250 22041
rect 5214 20619 5250 21251
rect 5214 19829 5250 20461
rect 5214 19039 5250 19671
rect 5214 18249 5250 18881
rect 5214 17459 5250 18091
rect 5214 16669 5250 17301
rect 5214 15879 5250 16511
rect 5214 15089 5250 15721
rect 5214 14299 5250 14931
rect 5214 13509 5250 14141
rect 5214 12719 5250 13351
rect 5214 11929 5250 12561
rect 5214 11139 5250 11771
rect 5214 10349 5250 10981
rect 5214 9559 5250 10191
rect 5214 8769 5250 9401
rect 5214 7979 5250 8611
rect 5214 7189 5250 7821
rect 5214 6399 5250 7031
rect 5214 5609 5250 6241
rect 5214 4819 5250 5451
rect 5214 4029 5250 4661
rect 5214 3239 5250 3871
rect 5214 2449 5250 3081
rect 5214 1659 5250 2291
rect 5214 869 5250 1501
rect 5214 79 5250 711
rect 5286 0 5322 25280
rect 5358 0 5394 25280
rect 5838 0 5874 25280
rect 5910 0 5946 25280
rect 5982 24569 6018 25201
rect 5982 23779 6018 24411
rect 5982 22989 6018 23621
rect 5982 22199 6018 22831
rect 5982 21409 6018 22041
rect 5982 20619 6018 21251
rect 5982 19829 6018 20461
rect 5982 19039 6018 19671
rect 5982 18249 6018 18881
rect 5982 17459 6018 18091
rect 5982 16669 6018 17301
rect 5982 15879 6018 16511
rect 5982 15089 6018 15721
rect 5982 14299 6018 14931
rect 5982 13509 6018 14141
rect 5982 12719 6018 13351
rect 5982 11929 6018 12561
rect 5982 11139 6018 11771
rect 5982 10349 6018 10981
rect 5982 9559 6018 10191
rect 5982 8769 6018 9401
rect 5982 7979 6018 8611
rect 5982 7189 6018 7821
rect 5982 6399 6018 7031
rect 5982 5609 6018 6241
rect 5982 4819 6018 5451
rect 5982 4029 6018 4661
rect 5982 3239 6018 3871
rect 5982 2449 6018 3081
rect 5982 1659 6018 2291
rect 5982 869 6018 1501
rect 5982 79 6018 711
rect 6054 0 6090 25280
rect 6126 0 6162 25280
rect 6318 0 6354 25280
rect 6390 0 6426 25280
rect 6462 24569 6498 25201
rect 6462 23779 6498 24411
rect 6462 22989 6498 23621
rect 6462 22199 6498 22831
rect 6462 21409 6498 22041
rect 6462 20619 6498 21251
rect 6462 19829 6498 20461
rect 6462 19039 6498 19671
rect 6462 18249 6498 18881
rect 6462 17459 6498 18091
rect 6462 16669 6498 17301
rect 6462 15879 6498 16511
rect 6462 15089 6498 15721
rect 6462 14299 6498 14931
rect 6462 13509 6498 14141
rect 6462 12719 6498 13351
rect 6462 11929 6498 12561
rect 6462 11139 6498 11771
rect 6462 10349 6498 10981
rect 6462 9559 6498 10191
rect 6462 8769 6498 9401
rect 6462 7979 6498 8611
rect 6462 7189 6498 7821
rect 6462 6399 6498 7031
rect 6462 5609 6498 6241
rect 6462 4819 6498 5451
rect 6462 4029 6498 4661
rect 6462 3239 6498 3871
rect 6462 2449 6498 3081
rect 6462 1659 6498 2291
rect 6462 869 6498 1501
rect 6462 79 6498 711
rect 6534 0 6570 25280
rect 6606 0 6642 25280
rect 7086 0 7122 25280
rect 7158 0 7194 25280
rect 7230 24569 7266 25201
rect 7230 23779 7266 24411
rect 7230 22989 7266 23621
rect 7230 22199 7266 22831
rect 7230 21409 7266 22041
rect 7230 20619 7266 21251
rect 7230 19829 7266 20461
rect 7230 19039 7266 19671
rect 7230 18249 7266 18881
rect 7230 17459 7266 18091
rect 7230 16669 7266 17301
rect 7230 15879 7266 16511
rect 7230 15089 7266 15721
rect 7230 14299 7266 14931
rect 7230 13509 7266 14141
rect 7230 12719 7266 13351
rect 7230 11929 7266 12561
rect 7230 11139 7266 11771
rect 7230 10349 7266 10981
rect 7230 9559 7266 10191
rect 7230 8769 7266 9401
rect 7230 7979 7266 8611
rect 7230 7189 7266 7821
rect 7230 6399 7266 7031
rect 7230 5609 7266 6241
rect 7230 4819 7266 5451
rect 7230 4029 7266 4661
rect 7230 3239 7266 3871
rect 7230 2449 7266 3081
rect 7230 1659 7266 2291
rect 7230 869 7266 1501
rect 7230 79 7266 711
rect 7302 0 7338 25280
rect 7374 0 7410 25280
rect 7566 0 7602 25280
rect 7638 0 7674 25280
rect 7710 24569 7746 25201
rect 7710 23779 7746 24411
rect 7710 22989 7746 23621
rect 7710 22199 7746 22831
rect 7710 21409 7746 22041
rect 7710 20619 7746 21251
rect 7710 19829 7746 20461
rect 7710 19039 7746 19671
rect 7710 18249 7746 18881
rect 7710 17459 7746 18091
rect 7710 16669 7746 17301
rect 7710 15879 7746 16511
rect 7710 15089 7746 15721
rect 7710 14299 7746 14931
rect 7710 13509 7746 14141
rect 7710 12719 7746 13351
rect 7710 11929 7746 12561
rect 7710 11139 7746 11771
rect 7710 10349 7746 10981
rect 7710 9559 7746 10191
rect 7710 8769 7746 9401
rect 7710 7979 7746 8611
rect 7710 7189 7746 7821
rect 7710 6399 7746 7031
rect 7710 5609 7746 6241
rect 7710 4819 7746 5451
rect 7710 4029 7746 4661
rect 7710 3239 7746 3871
rect 7710 2449 7746 3081
rect 7710 1659 7746 2291
rect 7710 869 7746 1501
rect 7710 79 7746 711
rect 7782 0 7818 25280
rect 7854 0 7890 25280
rect 8334 0 8370 25280
rect 8406 0 8442 25280
rect 8478 24569 8514 25201
rect 8478 23779 8514 24411
rect 8478 22989 8514 23621
rect 8478 22199 8514 22831
rect 8478 21409 8514 22041
rect 8478 20619 8514 21251
rect 8478 19829 8514 20461
rect 8478 19039 8514 19671
rect 8478 18249 8514 18881
rect 8478 17459 8514 18091
rect 8478 16669 8514 17301
rect 8478 15879 8514 16511
rect 8478 15089 8514 15721
rect 8478 14299 8514 14931
rect 8478 13509 8514 14141
rect 8478 12719 8514 13351
rect 8478 11929 8514 12561
rect 8478 11139 8514 11771
rect 8478 10349 8514 10981
rect 8478 9559 8514 10191
rect 8478 8769 8514 9401
rect 8478 7979 8514 8611
rect 8478 7189 8514 7821
rect 8478 6399 8514 7031
rect 8478 5609 8514 6241
rect 8478 4819 8514 5451
rect 8478 4029 8514 4661
rect 8478 3239 8514 3871
rect 8478 2449 8514 3081
rect 8478 1659 8514 2291
rect 8478 869 8514 1501
rect 8478 79 8514 711
rect 8550 0 8586 25280
rect 8622 0 8658 25280
rect 8814 0 8850 25280
rect 8886 0 8922 25280
rect 8958 24569 8994 25201
rect 8958 23779 8994 24411
rect 8958 22989 8994 23621
rect 8958 22199 8994 22831
rect 8958 21409 8994 22041
rect 8958 20619 8994 21251
rect 8958 19829 8994 20461
rect 8958 19039 8994 19671
rect 8958 18249 8994 18881
rect 8958 17459 8994 18091
rect 8958 16669 8994 17301
rect 8958 15879 8994 16511
rect 8958 15089 8994 15721
rect 8958 14299 8994 14931
rect 8958 13509 8994 14141
rect 8958 12719 8994 13351
rect 8958 11929 8994 12561
rect 8958 11139 8994 11771
rect 8958 10349 8994 10981
rect 8958 9559 8994 10191
rect 8958 8769 8994 9401
rect 8958 7979 8994 8611
rect 8958 7189 8994 7821
rect 8958 6399 8994 7031
rect 8958 5609 8994 6241
rect 8958 4819 8994 5451
rect 8958 4029 8994 4661
rect 8958 3239 8994 3871
rect 8958 2449 8994 3081
rect 8958 1659 8994 2291
rect 8958 869 8994 1501
rect 8958 79 8994 711
rect 9030 0 9066 25280
rect 9102 0 9138 25280
rect 9582 0 9618 25280
rect 9654 0 9690 25280
rect 9726 24569 9762 25201
rect 9726 23779 9762 24411
rect 9726 22989 9762 23621
rect 9726 22199 9762 22831
rect 9726 21409 9762 22041
rect 9726 20619 9762 21251
rect 9726 19829 9762 20461
rect 9726 19039 9762 19671
rect 9726 18249 9762 18881
rect 9726 17459 9762 18091
rect 9726 16669 9762 17301
rect 9726 15879 9762 16511
rect 9726 15089 9762 15721
rect 9726 14299 9762 14931
rect 9726 13509 9762 14141
rect 9726 12719 9762 13351
rect 9726 11929 9762 12561
rect 9726 11139 9762 11771
rect 9726 10349 9762 10981
rect 9726 9559 9762 10191
rect 9726 8769 9762 9401
rect 9726 7979 9762 8611
rect 9726 7189 9762 7821
rect 9726 6399 9762 7031
rect 9726 5609 9762 6241
rect 9726 4819 9762 5451
rect 9726 4029 9762 4661
rect 9726 3239 9762 3871
rect 9726 2449 9762 3081
rect 9726 1659 9762 2291
rect 9726 869 9762 1501
rect 9726 79 9762 711
rect 9798 0 9834 25280
rect 9870 0 9906 25280
rect 10062 0 10098 25280
rect 10134 0 10170 25280
rect 10206 24569 10242 25201
rect 10206 23779 10242 24411
rect 10206 22989 10242 23621
rect 10206 22199 10242 22831
rect 10206 21409 10242 22041
rect 10206 20619 10242 21251
rect 10206 19829 10242 20461
rect 10206 19039 10242 19671
rect 10206 18249 10242 18881
rect 10206 17459 10242 18091
rect 10206 16669 10242 17301
rect 10206 15879 10242 16511
rect 10206 15089 10242 15721
rect 10206 14299 10242 14931
rect 10206 13509 10242 14141
rect 10206 12719 10242 13351
rect 10206 11929 10242 12561
rect 10206 11139 10242 11771
rect 10206 10349 10242 10981
rect 10206 9559 10242 10191
rect 10206 8769 10242 9401
rect 10206 7979 10242 8611
rect 10206 7189 10242 7821
rect 10206 6399 10242 7031
rect 10206 5609 10242 6241
rect 10206 4819 10242 5451
rect 10206 4029 10242 4661
rect 10206 3239 10242 3871
rect 10206 2449 10242 3081
rect 10206 1659 10242 2291
rect 10206 869 10242 1501
rect 10206 79 10242 711
rect 10278 0 10314 25280
rect 10350 0 10386 25280
rect 10830 0 10866 25280
rect 10902 0 10938 25280
rect 10974 24569 11010 25201
rect 10974 23779 11010 24411
rect 10974 22989 11010 23621
rect 10974 22199 11010 22831
rect 10974 21409 11010 22041
rect 10974 20619 11010 21251
rect 10974 19829 11010 20461
rect 10974 19039 11010 19671
rect 10974 18249 11010 18881
rect 10974 17459 11010 18091
rect 10974 16669 11010 17301
rect 10974 15879 11010 16511
rect 10974 15089 11010 15721
rect 10974 14299 11010 14931
rect 10974 13509 11010 14141
rect 10974 12719 11010 13351
rect 10974 11929 11010 12561
rect 10974 11139 11010 11771
rect 10974 10349 11010 10981
rect 10974 9559 11010 10191
rect 10974 8769 11010 9401
rect 10974 7979 11010 8611
rect 10974 7189 11010 7821
rect 10974 6399 11010 7031
rect 10974 5609 11010 6241
rect 10974 4819 11010 5451
rect 10974 4029 11010 4661
rect 10974 3239 11010 3871
rect 10974 2449 11010 3081
rect 10974 1659 11010 2291
rect 10974 869 11010 1501
rect 10974 79 11010 711
rect 11046 0 11082 25280
rect 11118 0 11154 25280
rect 11310 0 11346 25280
rect 11382 0 11418 25280
rect 11454 24569 11490 25201
rect 11454 23779 11490 24411
rect 11454 22989 11490 23621
rect 11454 22199 11490 22831
rect 11454 21409 11490 22041
rect 11454 20619 11490 21251
rect 11454 19829 11490 20461
rect 11454 19039 11490 19671
rect 11454 18249 11490 18881
rect 11454 17459 11490 18091
rect 11454 16669 11490 17301
rect 11454 15879 11490 16511
rect 11454 15089 11490 15721
rect 11454 14299 11490 14931
rect 11454 13509 11490 14141
rect 11454 12719 11490 13351
rect 11454 11929 11490 12561
rect 11454 11139 11490 11771
rect 11454 10349 11490 10981
rect 11454 9559 11490 10191
rect 11454 8769 11490 9401
rect 11454 7979 11490 8611
rect 11454 7189 11490 7821
rect 11454 6399 11490 7031
rect 11454 5609 11490 6241
rect 11454 4819 11490 5451
rect 11454 4029 11490 4661
rect 11454 3239 11490 3871
rect 11454 2449 11490 3081
rect 11454 1659 11490 2291
rect 11454 869 11490 1501
rect 11454 79 11490 711
rect 11526 0 11562 25280
rect 11598 0 11634 25280
rect 12078 0 12114 25280
rect 12150 0 12186 25280
rect 12222 24569 12258 25201
rect 12222 23779 12258 24411
rect 12222 22989 12258 23621
rect 12222 22199 12258 22831
rect 12222 21409 12258 22041
rect 12222 20619 12258 21251
rect 12222 19829 12258 20461
rect 12222 19039 12258 19671
rect 12222 18249 12258 18881
rect 12222 17459 12258 18091
rect 12222 16669 12258 17301
rect 12222 15879 12258 16511
rect 12222 15089 12258 15721
rect 12222 14299 12258 14931
rect 12222 13509 12258 14141
rect 12222 12719 12258 13351
rect 12222 11929 12258 12561
rect 12222 11139 12258 11771
rect 12222 10349 12258 10981
rect 12222 9559 12258 10191
rect 12222 8769 12258 9401
rect 12222 7979 12258 8611
rect 12222 7189 12258 7821
rect 12222 6399 12258 7031
rect 12222 5609 12258 6241
rect 12222 4819 12258 5451
rect 12222 4029 12258 4661
rect 12222 3239 12258 3871
rect 12222 2449 12258 3081
rect 12222 1659 12258 2291
rect 12222 869 12258 1501
rect 12222 79 12258 711
rect 12294 0 12330 25280
rect 12366 0 12402 25280
rect 12558 0 12594 25280
rect 12630 0 12666 25280
rect 12702 24569 12738 25201
rect 12702 23779 12738 24411
rect 12702 22989 12738 23621
rect 12702 22199 12738 22831
rect 12702 21409 12738 22041
rect 12702 20619 12738 21251
rect 12702 19829 12738 20461
rect 12702 19039 12738 19671
rect 12702 18249 12738 18881
rect 12702 17459 12738 18091
rect 12702 16669 12738 17301
rect 12702 15879 12738 16511
rect 12702 15089 12738 15721
rect 12702 14299 12738 14931
rect 12702 13509 12738 14141
rect 12702 12719 12738 13351
rect 12702 11929 12738 12561
rect 12702 11139 12738 11771
rect 12702 10349 12738 10981
rect 12702 9559 12738 10191
rect 12702 8769 12738 9401
rect 12702 7979 12738 8611
rect 12702 7189 12738 7821
rect 12702 6399 12738 7031
rect 12702 5609 12738 6241
rect 12702 4819 12738 5451
rect 12702 4029 12738 4661
rect 12702 3239 12738 3871
rect 12702 2449 12738 3081
rect 12702 1659 12738 2291
rect 12702 869 12738 1501
rect 12702 79 12738 711
rect 12774 0 12810 25280
rect 12846 0 12882 25280
rect 13326 0 13362 25280
rect 13398 0 13434 25280
rect 13470 24569 13506 25201
rect 13470 23779 13506 24411
rect 13470 22989 13506 23621
rect 13470 22199 13506 22831
rect 13470 21409 13506 22041
rect 13470 20619 13506 21251
rect 13470 19829 13506 20461
rect 13470 19039 13506 19671
rect 13470 18249 13506 18881
rect 13470 17459 13506 18091
rect 13470 16669 13506 17301
rect 13470 15879 13506 16511
rect 13470 15089 13506 15721
rect 13470 14299 13506 14931
rect 13470 13509 13506 14141
rect 13470 12719 13506 13351
rect 13470 11929 13506 12561
rect 13470 11139 13506 11771
rect 13470 10349 13506 10981
rect 13470 9559 13506 10191
rect 13470 8769 13506 9401
rect 13470 7979 13506 8611
rect 13470 7189 13506 7821
rect 13470 6399 13506 7031
rect 13470 5609 13506 6241
rect 13470 4819 13506 5451
rect 13470 4029 13506 4661
rect 13470 3239 13506 3871
rect 13470 2449 13506 3081
rect 13470 1659 13506 2291
rect 13470 869 13506 1501
rect 13470 79 13506 711
rect 13542 0 13578 25280
rect 13614 0 13650 25280
rect 13806 0 13842 25280
rect 13878 0 13914 25280
rect 13950 24569 13986 25201
rect 13950 23779 13986 24411
rect 13950 22989 13986 23621
rect 13950 22199 13986 22831
rect 13950 21409 13986 22041
rect 13950 20619 13986 21251
rect 13950 19829 13986 20461
rect 13950 19039 13986 19671
rect 13950 18249 13986 18881
rect 13950 17459 13986 18091
rect 13950 16669 13986 17301
rect 13950 15879 13986 16511
rect 13950 15089 13986 15721
rect 13950 14299 13986 14931
rect 13950 13509 13986 14141
rect 13950 12719 13986 13351
rect 13950 11929 13986 12561
rect 13950 11139 13986 11771
rect 13950 10349 13986 10981
rect 13950 9559 13986 10191
rect 13950 8769 13986 9401
rect 13950 7979 13986 8611
rect 13950 7189 13986 7821
rect 13950 6399 13986 7031
rect 13950 5609 13986 6241
rect 13950 4819 13986 5451
rect 13950 4029 13986 4661
rect 13950 3239 13986 3871
rect 13950 2449 13986 3081
rect 13950 1659 13986 2291
rect 13950 869 13986 1501
rect 13950 79 13986 711
rect 14022 0 14058 25280
rect 14094 0 14130 25280
rect 14574 0 14610 25280
rect 14646 0 14682 25280
rect 14718 24569 14754 25201
rect 14718 23779 14754 24411
rect 14718 22989 14754 23621
rect 14718 22199 14754 22831
rect 14718 21409 14754 22041
rect 14718 20619 14754 21251
rect 14718 19829 14754 20461
rect 14718 19039 14754 19671
rect 14718 18249 14754 18881
rect 14718 17459 14754 18091
rect 14718 16669 14754 17301
rect 14718 15879 14754 16511
rect 14718 15089 14754 15721
rect 14718 14299 14754 14931
rect 14718 13509 14754 14141
rect 14718 12719 14754 13351
rect 14718 11929 14754 12561
rect 14718 11139 14754 11771
rect 14718 10349 14754 10981
rect 14718 9559 14754 10191
rect 14718 8769 14754 9401
rect 14718 7979 14754 8611
rect 14718 7189 14754 7821
rect 14718 6399 14754 7031
rect 14718 5609 14754 6241
rect 14718 4819 14754 5451
rect 14718 4029 14754 4661
rect 14718 3239 14754 3871
rect 14718 2449 14754 3081
rect 14718 1659 14754 2291
rect 14718 869 14754 1501
rect 14718 79 14754 711
rect 14790 0 14826 25280
rect 14862 0 14898 25280
rect 15054 0 15090 25280
rect 15126 0 15162 25280
rect 15198 24569 15234 25201
rect 15198 23779 15234 24411
rect 15198 22989 15234 23621
rect 15198 22199 15234 22831
rect 15198 21409 15234 22041
rect 15198 20619 15234 21251
rect 15198 19829 15234 20461
rect 15198 19039 15234 19671
rect 15198 18249 15234 18881
rect 15198 17459 15234 18091
rect 15198 16669 15234 17301
rect 15198 15879 15234 16511
rect 15198 15089 15234 15721
rect 15198 14299 15234 14931
rect 15198 13509 15234 14141
rect 15198 12719 15234 13351
rect 15198 11929 15234 12561
rect 15198 11139 15234 11771
rect 15198 10349 15234 10981
rect 15198 9559 15234 10191
rect 15198 8769 15234 9401
rect 15198 7979 15234 8611
rect 15198 7189 15234 7821
rect 15198 6399 15234 7031
rect 15198 5609 15234 6241
rect 15198 4819 15234 5451
rect 15198 4029 15234 4661
rect 15198 3239 15234 3871
rect 15198 2449 15234 3081
rect 15198 1659 15234 2291
rect 15198 869 15234 1501
rect 15198 79 15234 711
rect 15270 0 15306 25280
rect 15342 0 15378 25280
rect 15822 0 15858 25280
rect 15894 0 15930 25280
rect 15966 24569 16002 25201
rect 15966 23779 16002 24411
rect 15966 22989 16002 23621
rect 15966 22199 16002 22831
rect 15966 21409 16002 22041
rect 15966 20619 16002 21251
rect 15966 19829 16002 20461
rect 15966 19039 16002 19671
rect 15966 18249 16002 18881
rect 15966 17459 16002 18091
rect 15966 16669 16002 17301
rect 15966 15879 16002 16511
rect 15966 15089 16002 15721
rect 15966 14299 16002 14931
rect 15966 13509 16002 14141
rect 15966 12719 16002 13351
rect 15966 11929 16002 12561
rect 15966 11139 16002 11771
rect 15966 10349 16002 10981
rect 15966 9559 16002 10191
rect 15966 8769 16002 9401
rect 15966 7979 16002 8611
rect 15966 7189 16002 7821
rect 15966 6399 16002 7031
rect 15966 5609 16002 6241
rect 15966 4819 16002 5451
rect 15966 4029 16002 4661
rect 15966 3239 16002 3871
rect 15966 2449 16002 3081
rect 15966 1659 16002 2291
rect 15966 869 16002 1501
rect 15966 79 16002 711
rect 16038 0 16074 25280
rect 16110 0 16146 25280
rect 16302 0 16338 25280
rect 16374 0 16410 25280
rect 16446 24569 16482 25201
rect 16446 23779 16482 24411
rect 16446 22989 16482 23621
rect 16446 22199 16482 22831
rect 16446 21409 16482 22041
rect 16446 20619 16482 21251
rect 16446 19829 16482 20461
rect 16446 19039 16482 19671
rect 16446 18249 16482 18881
rect 16446 17459 16482 18091
rect 16446 16669 16482 17301
rect 16446 15879 16482 16511
rect 16446 15089 16482 15721
rect 16446 14299 16482 14931
rect 16446 13509 16482 14141
rect 16446 12719 16482 13351
rect 16446 11929 16482 12561
rect 16446 11139 16482 11771
rect 16446 10349 16482 10981
rect 16446 9559 16482 10191
rect 16446 8769 16482 9401
rect 16446 7979 16482 8611
rect 16446 7189 16482 7821
rect 16446 6399 16482 7031
rect 16446 5609 16482 6241
rect 16446 4819 16482 5451
rect 16446 4029 16482 4661
rect 16446 3239 16482 3871
rect 16446 2449 16482 3081
rect 16446 1659 16482 2291
rect 16446 869 16482 1501
rect 16446 79 16482 711
rect 16518 0 16554 25280
rect 16590 0 16626 25280
rect 17070 0 17106 25280
rect 17142 0 17178 25280
rect 17214 24569 17250 25201
rect 17214 23779 17250 24411
rect 17214 22989 17250 23621
rect 17214 22199 17250 22831
rect 17214 21409 17250 22041
rect 17214 20619 17250 21251
rect 17214 19829 17250 20461
rect 17214 19039 17250 19671
rect 17214 18249 17250 18881
rect 17214 17459 17250 18091
rect 17214 16669 17250 17301
rect 17214 15879 17250 16511
rect 17214 15089 17250 15721
rect 17214 14299 17250 14931
rect 17214 13509 17250 14141
rect 17214 12719 17250 13351
rect 17214 11929 17250 12561
rect 17214 11139 17250 11771
rect 17214 10349 17250 10981
rect 17214 9559 17250 10191
rect 17214 8769 17250 9401
rect 17214 7979 17250 8611
rect 17214 7189 17250 7821
rect 17214 6399 17250 7031
rect 17214 5609 17250 6241
rect 17214 4819 17250 5451
rect 17214 4029 17250 4661
rect 17214 3239 17250 3871
rect 17214 2449 17250 3081
rect 17214 1659 17250 2291
rect 17214 869 17250 1501
rect 17214 79 17250 711
rect 17286 0 17322 25280
rect 17358 0 17394 25280
rect 17550 0 17586 25280
rect 17622 0 17658 25280
rect 17694 24569 17730 25201
rect 17694 23779 17730 24411
rect 17694 22989 17730 23621
rect 17694 22199 17730 22831
rect 17694 21409 17730 22041
rect 17694 20619 17730 21251
rect 17694 19829 17730 20461
rect 17694 19039 17730 19671
rect 17694 18249 17730 18881
rect 17694 17459 17730 18091
rect 17694 16669 17730 17301
rect 17694 15879 17730 16511
rect 17694 15089 17730 15721
rect 17694 14299 17730 14931
rect 17694 13509 17730 14141
rect 17694 12719 17730 13351
rect 17694 11929 17730 12561
rect 17694 11139 17730 11771
rect 17694 10349 17730 10981
rect 17694 9559 17730 10191
rect 17694 8769 17730 9401
rect 17694 7979 17730 8611
rect 17694 7189 17730 7821
rect 17694 6399 17730 7031
rect 17694 5609 17730 6241
rect 17694 4819 17730 5451
rect 17694 4029 17730 4661
rect 17694 3239 17730 3871
rect 17694 2449 17730 3081
rect 17694 1659 17730 2291
rect 17694 869 17730 1501
rect 17694 79 17730 711
rect 17766 0 17802 25280
rect 17838 0 17874 25280
rect 18318 0 18354 25280
rect 18390 0 18426 25280
rect 18462 24569 18498 25201
rect 18462 23779 18498 24411
rect 18462 22989 18498 23621
rect 18462 22199 18498 22831
rect 18462 21409 18498 22041
rect 18462 20619 18498 21251
rect 18462 19829 18498 20461
rect 18462 19039 18498 19671
rect 18462 18249 18498 18881
rect 18462 17459 18498 18091
rect 18462 16669 18498 17301
rect 18462 15879 18498 16511
rect 18462 15089 18498 15721
rect 18462 14299 18498 14931
rect 18462 13509 18498 14141
rect 18462 12719 18498 13351
rect 18462 11929 18498 12561
rect 18462 11139 18498 11771
rect 18462 10349 18498 10981
rect 18462 9559 18498 10191
rect 18462 8769 18498 9401
rect 18462 7979 18498 8611
rect 18462 7189 18498 7821
rect 18462 6399 18498 7031
rect 18462 5609 18498 6241
rect 18462 4819 18498 5451
rect 18462 4029 18498 4661
rect 18462 3239 18498 3871
rect 18462 2449 18498 3081
rect 18462 1659 18498 2291
rect 18462 869 18498 1501
rect 18462 79 18498 711
rect 18534 0 18570 25280
rect 18606 0 18642 25280
rect 18798 0 18834 25280
rect 18870 0 18906 25280
rect 18942 24569 18978 25201
rect 18942 23779 18978 24411
rect 18942 22989 18978 23621
rect 18942 22199 18978 22831
rect 18942 21409 18978 22041
rect 18942 20619 18978 21251
rect 18942 19829 18978 20461
rect 18942 19039 18978 19671
rect 18942 18249 18978 18881
rect 18942 17459 18978 18091
rect 18942 16669 18978 17301
rect 18942 15879 18978 16511
rect 18942 15089 18978 15721
rect 18942 14299 18978 14931
rect 18942 13509 18978 14141
rect 18942 12719 18978 13351
rect 18942 11929 18978 12561
rect 18942 11139 18978 11771
rect 18942 10349 18978 10981
rect 18942 9559 18978 10191
rect 18942 8769 18978 9401
rect 18942 7979 18978 8611
rect 18942 7189 18978 7821
rect 18942 6399 18978 7031
rect 18942 5609 18978 6241
rect 18942 4819 18978 5451
rect 18942 4029 18978 4661
rect 18942 3239 18978 3871
rect 18942 2449 18978 3081
rect 18942 1659 18978 2291
rect 18942 869 18978 1501
rect 18942 79 18978 711
rect 19014 0 19050 25280
rect 19086 0 19122 25280
rect 19566 0 19602 25280
rect 19638 0 19674 25280
rect 19710 24569 19746 25201
rect 19710 23779 19746 24411
rect 19710 22989 19746 23621
rect 19710 22199 19746 22831
rect 19710 21409 19746 22041
rect 19710 20619 19746 21251
rect 19710 19829 19746 20461
rect 19710 19039 19746 19671
rect 19710 18249 19746 18881
rect 19710 17459 19746 18091
rect 19710 16669 19746 17301
rect 19710 15879 19746 16511
rect 19710 15089 19746 15721
rect 19710 14299 19746 14931
rect 19710 13509 19746 14141
rect 19710 12719 19746 13351
rect 19710 11929 19746 12561
rect 19710 11139 19746 11771
rect 19710 10349 19746 10981
rect 19710 9559 19746 10191
rect 19710 8769 19746 9401
rect 19710 7979 19746 8611
rect 19710 7189 19746 7821
rect 19710 6399 19746 7031
rect 19710 5609 19746 6241
rect 19710 4819 19746 5451
rect 19710 4029 19746 4661
rect 19710 3239 19746 3871
rect 19710 2449 19746 3081
rect 19710 1659 19746 2291
rect 19710 869 19746 1501
rect 19710 79 19746 711
rect 19782 0 19818 25280
rect 19854 0 19890 25280
<< metal2 >>
rect 186 25225 294 25335
rect 954 25225 1062 25335
rect 1434 25225 1542 25335
rect 2202 25225 2310 25335
rect 2682 25225 2790 25335
rect 3450 25225 3558 25335
rect 3930 25225 4038 25335
rect 4698 25225 4806 25335
rect 5178 25225 5286 25335
rect 5946 25225 6054 25335
rect 6426 25225 6534 25335
rect 7194 25225 7302 25335
rect 7674 25225 7782 25335
rect 8442 25225 8550 25335
rect 8922 25225 9030 25335
rect 9690 25225 9798 25335
rect 10170 25225 10278 25335
rect 10938 25225 11046 25335
rect 11418 25225 11526 25335
rect 12186 25225 12294 25335
rect 12666 25225 12774 25335
rect 13434 25225 13542 25335
rect 13914 25225 14022 25335
rect 14682 25225 14790 25335
rect 15162 25225 15270 25335
rect 15930 25225 16038 25335
rect 16410 25225 16518 25335
rect 17178 25225 17286 25335
rect 17658 25225 17766 25335
rect 18426 25225 18534 25335
rect 18906 25225 19014 25335
rect 19674 25225 19782 25335
rect 0 25129 19968 25177
rect 186 25005 294 25081
rect 954 25005 1062 25081
rect 1434 25005 1542 25081
rect 2202 25005 2310 25081
rect 2682 25005 2790 25081
rect 3450 25005 3558 25081
rect 3930 25005 4038 25081
rect 4698 25005 4806 25081
rect 5178 25005 5286 25081
rect 5946 25005 6054 25081
rect 6426 25005 6534 25081
rect 7194 25005 7302 25081
rect 7674 25005 7782 25081
rect 8442 25005 8550 25081
rect 8922 25005 9030 25081
rect 9690 25005 9798 25081
rect 10170 25005 10278 25081
rect 10938 25005 11046 25081
rect 11418 25005 11526 25081
rect 12186 25005 12294 25081
rect 12666 25005 12774 25081
rect 13434 25005 13542 25081
rect 13914 25005 14022 25081
rect 14682 25005 14790 25081
rect 15162 25005 15270 25081
rect 15930 25005 16038 25081
rect 16410 25005 16518 25081
rect 17178 25005 17286 25081
rect 17658 25005 17766 25081
rect 18426 25005 18534 25081
rect 18906 25005 19014 25081
rect 19674 25005 19782 25081
rect 0 24909 19968 24957
rect 0 24813 19968 24861
rect 186 24689 294 24765
rect 954 24689 1062 24765
rect 1434 24689 1542 24765
rect 2202 24689 2310 24765
rect 2682 24689 2790 24765
rect 3450 24689 3558 24765
rect 3930 24689 4038 24765
rect 4698 24689 4806 24765
rect 5178 24689 5286 24765
rect 5946 24689 6054 24765
rect 6426 24689 6534 24765
rect 7194 24689 7302 24765
rect 7674 24689 7782 24765
rect 8442 24689 8550 24765
rect 8922 24689 9030 24765
rect 9690 24689 9798 24765
rect 10170 24689 10278 24765
rect 10938 24689 11046 24765
rect 11418 24689 11526 24765
rect 12186 24689 12294 24765
rect 12666 24689 12774 24765
rect 13434 24689 13542 24765
rect 13914 24689 14022 24765
rect 14682 24689 14790 24765
rect 15162 24689 15270 24765
rect 15930 24689 16038 24765
rect 16410 24689 16518 24765
rect 17178 24689 17286 24765
rect 17658 24689 17766 24765
rect 18426 24689 18534 24765
rect 18906 24689 19014 24765
rect 19674 24689 19782 24765
rect 0 24593 19968 24641
rect 186 24435 294 24545
rect 954 24435 1062 24545
rect 1434 24435 1542 24545
rect 2202 24435 2310 24545
rect 2682 24435 2790 24545
rect 3450 24435 3558 24545
rect 3930 24435 4038 24545
rect 4698 24435 4806 24545
rect 5178 24435 5286 24545
rect 5946 24435 6054 24545
rect 6426 24435 6534 24545
rect 7194 24435 7302 24545
rect 7674 24435 7782 24545
rect 8442 24435 8550 24545
rect 8922 24435 9030 24545
rect 9690 24435 9798 24545
rect 10170 24435 10278 24545
rect 10938 24435 11046 24545
rect 11418 24435 11526 24545
rect 12186 24435 12294 24545
rect 12666 24435 12774 24545
rect 13434 24435 13542 24545
rect 13914 24435 14022 24545
rect 14682 24435 14790 24545
rect 15162 24435 15270 24545
rect 15930 24435 16038 24545
rect 16410 24435 16518 24545
rect 17178 24435 17286 24545
rect 17658 24435 17766 24545
rect 18426 24435 18534 24545
rect 18906 24435 19014 24545
rect 19674 24435 19782 24545
rect 0 24339 19968 24387
rect 186 24215 294 24291
rect 954 24215 1062 24291
rect 1434 24215 1542 24291
rect 2202 24215 2310 24291
rect 2682 24215 2790 24291
rect 3450 24215 3558 24291
rect 3930 24215 4038 24291
rect 4698 24215 4806 24291
rect 5178 24215 5286 24291
rect 5946 24215 6054 24291
rect 6426 24215 6534 24291
rect 7194 24215 7302 24291
rect 7674 24215 7782 24291
rect 8442 24215 8550 24291
rect 8922 24215 9030 24291
rect 9690 24215 9798 24291
rect 10170 24215 10278 24291
rect 10938 24215 11046 24291
rect 11418 24215 11526 24291
rect 12186 24215 12294 24291
rect 12666 24215 12774 24291
rect 13434 24215 13542 24291
rect 13914 24215 14022 24291
rect 14682 24215 14790 24291
rect 15162 24215 15270 24291
rect 15930 24215 16038 24291
rect 16410 24215 16518 24291
rect 17178 24215 17286 24291
rect 17658 24215 17766 24291
rect 18426 24215 18534 24291
rect 18906 24215 19014 24291
rect 19674 24215 19782 24291
rect 0 24119 19968 24167
rect 0 24023 19968 24071
rect 186 23899 294 23975
rect 954 23899 1062 23975
rect 1434 23899 1542 23975
rect 2202 23899 2310 23975
rect 2682 23899 2790 23975
rect 3450 23899 3558 23975
rect 3930 23899 4038 23975
rect 4698 23899 4806 23975
rect 5178 23899 5286 23975
rect 5946 23899 6054 23975
rect 6426 23899 6534 23975
rect 7194 23899 7302 23975
rect 7674 23899 7782 23975
rect 8442 23899 8550 23975
rect 8922 23899 9030 23975
rect 9690 23899 9798 23975
rect 10170 23899 10278 23975
rect 10938 23899 11046 23975
rect 11418 23899 11526 23975
rect 12186 23899 12294 23975
rect 12666 23899 12774 23975
rect 13434 23899 13542 23975
rect 13914 23899 14022 23975
rect 14682 23899 14790 23975
rect 15162 23899 15270 23975
rect 15930 23899 16038 23975
rect 16410 23899 16518 23975
rect 17178 23899 17286 23975
rect 17658 23899 17766 23975
rect 18426 23899 18534 23975
rect 18906 23899 19014 23975
rect 19674 23899 19782 23975
rect 0 23803 19968 23851
rect 186 23645 294 23755
rect 954 23645 1062 23755
rect 1434 23645 1542 23755
rect 2202 23645 2310 23755
rect 2682 23645 2790 23755
rect 3450 23645 3558 23755
rect 3930 23645 4038 23755
rect 4698 23645 4806 23755
rect 5178 23645 5286 23755
rect 5946 23645 6054 23755
rect 6426 23645 6534 23755
rect 7194 23645 7302 23755
rect 7674 23645 7782 23755
rect 8442 23645 8550 23755
rect 8922 23645 9030 23755
rect 9690 23645 9798 23755
rect 10170 23645 10278 23755
rect 10938 23645 11046 23755
rect 11418 23645 11526 23755
rect 12186 23645 12294 23755
rect 12666 23645 12774 23755
rect 13434 23645 13542 23755
rect 13914 23645 14022 23755
rect 14682 23645 14790 23755
rect 15162 23645 15270 23755
rect 15930 23645 16038 23755
rect 16410 23645 16518 23755
rect 17178 23645 17286 23755
rect 17658 23645 17766 23755
rect 18426 23645 18534 23755
rect 18906 23645 19014 23755
rect 19674 23645 19782 23755
rect 0 23549 19968 23597
rect 186 23425 294 23501
rect 954 23425 1062 23501
rect 1434 23425 1542 23501
rect 2202 23425 2310 23501
rect 2682 23425 2790 23501
rect 3450 23425 3558 23501
rect 3930 23425 4038 23501
rect 4698 23425 4806 23501
rect 5178 23425 5286 23501
rect 5946 23425 6054 23501
rect 6426 23425 6534 23501
rect 7194 23425 7302 23501
rect 7674 23425 7782 23501
rect 8442 23425 8550 23501
rect 8922 23425 9030 23501
rect 9690 23425 9798 23501
rect 10170 23425 10278 23501
rect 10938 23425 11046 23501
rect 11418 23425 11526 23501
rect 12186 23425 12294 23501
rect 12666 23425 12774 23501
rect 13434 23425 13542 23501
rect 13914 23425 14022 23501
rect 14682 23425 14790 23501
rect 15162 23425 15270 23501
rect 15930 23425 16038 23501
rect 16410 23425 16518 23501
rect 17178 23425 17286 23501
rect 17658 23425 17766 23501
rect 18426 23425 18534 23501
rect 18906 23425 19014 23501
rect 19674 23425 19782 23501
rect 0 23329 19968 23377
rect 0 23233 19968 23281
rect 186 23109 294 23185
rect 954 23109 1062 23185
rect 1434 23109 1542 23185
rect 2202 23109 2310 23185
rect 2682 23109 2790 23185
rect 3450 23109 3558 23185
rect 3930 23109 4038 23185
rect 4698 23109 4806 23185
rect 5178 23109 5286 23185
rect 5946 23109 6054 23185
rect 6426 23109 6534 23185
rect 7194 23109 7302 23185
rect 7674 23109 7782 23185
rect 8442 23109 8550 23185
rect 8922 23109 9030 23185
rect 9690 23109 9798 23185
rect 10170 23109 10278 23185
rect 10938 23109 11046 23185
rect 11418 23109 11526 23185
rect 12186 23109 12294 23185
rect 12666 23109 12774 23185
rect 13434 23109 13542 23185
rect 13914 23109 14022 23185
rect 14682 23109 14790 23185
rect 15162 23109 15270 23185
rect 15930 23109 16038 23185
rect 16410 23109 16518 23185
rect 17178 23109 17286 23185
rect 17658 23109 17766 23185
rect 18426 23109 18534 23185
rect 18906 23109 19014 23185
rect 19674 23109 19782 23185
rect 0 23013 19968 23061
rect 186 22855 294 22965
rect 954 22855 1062 22965
rect 1434 22855 1542 22965
rect 2202 22855 2310 22965
rect 2682 22855 2790 22965
rect 3450 22855 3558 22965
rect 3930 22855 4038 22965
rect 4698 22855 4806 22965
rect 5178 22855 5286 22965
rect 5946 22855 6054 22965
rect 6426 22855 6534 22965
rect 7194 22855 7302 22965
rect 7674 22855 7782 22965
rect 8442 22855 8550 22965
rect 8922 22855 9030 22965
rect 9690 22855 9798 22965
rect 10170 22855 10278 22965
rect 10938 22855 11046 22965
rect 11418 22855 11526 22965
rect 12186 22855 12294 22965
rect 12666 22855 12774 22965
rect 13434 22855 13542 22965
rect 13914 22855 14022 22965
rect 14682 22855 14790 22965
rect 15162 22855 15270 22965
rect 15930 22855 16038 22965
rect 16410 22855 16518 22965
rect 17178 22855 17286 22965
rect 17658 22855 17766 22965
rect 18426 22855 18534 22965
rect 18906 22855 19014 22965
rect 19674 22855 19782 22965
rect 0 22759 19968 22807
rect 186 22635 294 22711
rect 954 22635 1062 22711
rect 1434 22635 1542 22711
rect 2202 22635 2310 22711
rect 2682 22635 2790 22711
rect 3450 22635 3558 22711
rect 3930 22635 4038 22711
rect 4698 22635 4806 22711
rect 5178 22635 5286 22711
rect 5946 22635 6054 22711
rect 6426 22635 6534 22711
rect 7194 22635 7302 22711
rect 7674 22635 7782 22711
rect 8442 22635 8550 22711
rect 8922 22635 9030 22711
rect 9690 22635 9798 22711
rect 10170 22635 10278 22711
rect 10938 22635 11046 22711
rect 11418 22635 11526 22711
rect 12186 22635 12294 22711
rect 12666 22635 12774 22711
rect 13434 22635 13542 22711
rect 13914 22635 14022 22711
rect 14682 22635 14790 22711
rect 15162 22635 15270 22711
rect 15930 22635 16038 22711
rect 16410 22635 16518 22711
rect 17178 22635 17286 22711
rect 17658 22635 17766 22711
rect 18426 22635 18534 22711
rect 18906 22635 19014 22711
rect 19674 22635 19782 22711
rect 0 22539 19968 22587
rect 0 22443 19968 22491
rect 186 22319 294 22395
rect 954 22319 1062 22395
rect 1434 22319 1542 22395
rect 2202 22319 2310 22395
rect 2682 22319 2790 22395
rect 3450 22319 3558 22395
rect 3930 22319 4038 22395
rect 4698 22319 4806 22395
rect 5178 22319 5286 22395
rect 5946 22319 6054 22395
rect 6426 22319 6534 22395
rect 7194 22319 7302 22395
rect 7674 22319 7782 22395
rect 8442 22319 8550 22395
rect 8922 22319 9030 22395
rect 9690 22319 9798 22395
rect 10170 22319 10278 22395
rect 10938 22319 11046 22395
rect 11418 22319 11526 22395
rect 12186 22319 12294 22395
rect 12666 22319 12774 22395
rect 13434 22319 13542 22395
rect 13914 22319 14022 22395
rect 14682 22319 14790 22395
rect 15162 22319 15270 22395
rect 15930 22319 16038 22395
rect 16410 22319 16518 22395
rect 17178 22319 17286 22395
rect 17658 22319 17766 22395
rect 18426 22319 18534 22395
rect 18906 22319 19014 22395
rect 19674 22319 19782 22395
rect 0 22223 19968 22271
rect 186 22065 294 22175
rect 954 22065 1062 22175
rect 1434 22065 1542 22175
rect 2202 22065 2310 22175
rect 2682 22065 2790 22175
rect 3450 22065 3558 22175
rect 3930 22065 4038 22175
rect 4698 22065 4806 22175
rect 5178 22065 5286 22175
rect 5946 22065 6054 22175
rect 6426 22065 6534 22175
rect 7194 22065 7302 22175
rect 7674 22065 7782 22175
rect 8442 22065 8550 22175
rect 8922 22065 9030 22175
rect 9690 22065 9798 22175
rect 10170 22065 10278 22175
rect 10938 22065 11046 22175
rect 11418 22065 11526 22175
rect 12186 22065 12294 22175
rect 12666 22065 12774 22175
rect 13434 22065 13542 22175
rect 13914 22065 14022 22175
rect 14682 22065 14790 22175
rect 15162 22065 15270 22175
rect 15930 22065 16038 22175
rect 16410 22065 16518 22175
rect 17178 22065 17286 22175
rect 17658 22065 17766 22175
rect 18426 22065 18534 22175
rect 18906 22065 19014 22175
rect 19674 22065 19782 22175
rect 0 21969 19968 22017
rect 186 21845 294 21921
rect 954 21845 1062 21921
rect 1434 21845 1542 21921
rect 2202 21845 2310 21921
rect 2682 21845 2790 21921
rect 3450 21845 3558 21921
rect 3930 21845 4038 21921
rect 4698 21845 4806 21921
rect 5178 21845 5286 21921
rect 5946 21845 6054 21921
rect 6426 21845 6534 21921
rect 7194 21845 7302 21921
rect 7674 21845 7782 21921
rect 8442 21845 8550 21921
rect 8922 21845 9030 21921
rect 9690 21845 9798 21921
rect 10170 21845 10278 21921
rect 10938 21845 11046 21921
rect 11418 21845 11526 21921
rect 12186 21845 12294 21921
rect 12666 21845 12774 21921
rect 13434 21845 13542 21921
rect 13914 21845 14022 21921
rect 14682 21845 14790 21921
rect 15162 21845 15270 21921
rect 15930 21845 16038 21921
rect 16410 21845 16518 21921
rect 17178 21845 17286 21921
rect 17658 21845 17766 21921
rect 18426 21845 18534 21921
rect 18906 21845 19014 21921
rect 19674 21845 19782 21921
rect 0 21749 19968 21797
rect 0 21653 19968 21701
rect 186 21529 294 21605
rect 954 21529 1062 21605
rect 1434 21529 1542 21605
rect 2202 21529 2310 21605
rect 2682 21529 2790 21605
rect 3450 21529 3558 21605
rect 3930 21529 4038 21605
rect 4698 21529 4806 21605
rect 5178 21529 5286 21605
rect 5946 21529 6054 21605
rect 6426 21529 6534 21605
rect 7194 21529 7302 21605
rect 7674 21529 7782 21605
rect 8442 21529 8550 21605
rect 8922 21529 9030 21605
rect 9690 21529 9798 21605
rect 10170 21529 10278 21605
rect 10938 21529 11046 21605
rect 11418 21529 11526 21605
rect 12186 21529 12294 21605
rect 12666 21529 12774 21605
rect 13434 21529 13542 21605
rect 13914 21529 14022 21605
rect 14682 21529 14790 21605
rect 15162 21529 15270 21605
rect 15930 21529 16038 21605
rect 16410 21529 16518 21605
rect 17178 21529 17286 21605
rect 17658 21529 17766 21605
rect 18426 21529 18534 21605
rect 18906 21529 19014 21605
rect 19674 21529 19782 21605
rect 0 21433 19968 21481
rect 186 21275 294 21385
rect 954 21275 1062 21385
rect 1434 21275 1542 21385
rect 2202 21275 2310 21385
rect 2682 21275 2790 21385
rect 3450 21275 3558 21385
rect 3930 21275 4038 21385
rect 4698 21275 4806 21385
rect 5178 21275 5286 21385
rect 5946 21275 6054 21385
rect 6426 21275 6534 21385
rect 7194 21275 7302 21385
rect 7674 21275 7782 21385
rect 8442 21275 8550 21385
rect 8922 21275 9030 21385
rect 9690 21275 9798 21385
rect 10170 21275 10278 21385
rect 10938 21275 11046 21385
rect 11418 21275 11526 21385
rect 12186 21275 12294 21385
rect 12666 21275 12774 21385
rect 13434 21275 13542 21385
rect 13914 21275 14022 21385
rect 14682 21275 14790 21385
rect 15162 21275 15270 21385
rect 15930 21275 16038 21385
rect 16410 21275 16518 21385
rect 17178 21275 17286 21385
rect 17658 21275 17766 21385
rect 18426 21275 18534 21385
rect 18906 21275 19014 21385
rect 19674 21275 19782 21385
rect 0 21179 19968 21227
rect 186 21055 294 21131
rect 954 21055 1062 21131
rect 1434 21055 1542 21131
rect 2202 21055 2310 21131
rect 2682 21055 2790 21131
rect 3450 21055 3558 21131
rect 3930 21055 4038 21131
rect 4698 21055 4806 21131
rect 5178 21055 5286 21131
rect 5946 21055 6054 21131
rect 6426 21055 6534 21131
rect 7194 21055 7302 21131
rect 7674 21055 7782 21131
rect 8442 21055 8550 21131
rect 8922 21055 9030 21131
rect 9690 21055 9798 21131
rect 10170 21055 10278 21131
rect 10938 21055 11046 21131
rect 11418 21055 11526 21131
rect 12186 21055 12294 21131
rect 12666 21055 12774 21131
rect 13434 21055 13542 21131
rect 13914 21055 14022 21131
rect 14682 21055 14790 21131
rect 15162 21055 15270 21131
rect 15930 21055 16038 21131
rect 16410 21055 16518 21131
rect 17178 21055 17286 21131
rect 17658 21055 17766 21131
rect 18426 21055 18534 21131
rect 18906 21055 19014 21131
rect 19674 21055 19782 21131
rect 0 20959 19968 21007
rect 0 20863 19968 20911
rect 186 20739 294 20815
rect 954 20739 1062 20815
rect 1434 20739 1542 20815
rect 2202 20739 2310 20815
rect 2682 20739 2790 20815
rect 3450 20739 3558 20815
rect 3930 20739 4038 20815
rect 4698 20739 4806 20815
rect 5178 20739 5286 20815
rect 5946 20739 6054 20815
rect 6426 20739 6534 20815
rect 7194 20739 7302 20815
rect 7674 20739 7782 20815
rect 8442 20739 8550 20815
rect 8922 20739 9030 20815
rect 9690 20739 9798 20815
rect 10170 20739 10278 20815
rect 10938 20739 11046 20815
rect 11418 20739 11526 20815
rect 12186 20739 12294 20815
rect 12666 20739 12774 20815
rect 13434 20739 13542 20815
rect 13914 20739 14022 20815
rect 14682 20739 14790 20815
rect 15162 20739 15270 20815
rect 15930 20739 16038 20815
rect 16410 20739 16518 20815
rect 17178 20739 17286 20815
rect 17658 20739 17766 20815
rect 18426 20739 18534 20815
rect 18906 20739 19014 20815
rect 19674 20739 19782 20815
rect 0 20643 19968 20691
rect 186 20485 294 20595
rect 954 20485 1062 20595
rect 1434 20485 1542 20595
rect 2202 20485 2310 20595
rect 2682 20485 2790 20595
rect 3450 20485 3558 20595
rect 3930 20485 4038 20595
rect 4698 20485 4806 20595
rect 5178 20485 5286 20595
rect 5946 20485 6054 20595
rect 6426 20485 6534 20595
rect 7194 20485 7302 20595
rect 7674 20485 7782 20595
rect 8442 20485 8550 20595
rect 8922 20485 9030 20595
rect 9690 20485 9798 20595
rect 10170 20485 10278 20595
rect 10938 20485 11046 20595
rect 11418 20485 11526 20595
rect 12186 20485 12294 20595
rect 12666 20485 12774 20595
rect 13434 20485 13542 20595
rect 13914 20485 14022 20595
rect 14682 20485 14790 20595
rect 15162 20485 15270 20595
rect 15930 20485 16038 20595
rect 16410 20485 16518 20595
rect 17178 20485 17286 20595
rect 17658 20485 17766 20595
rect 18426 20485 18534 20595
rect 18906 20485 19014 20595
rect 19674 20485 19782 20595
rect 0 20389 19968 20437
rect 186 20265 294 20341
rect 954 20265 1062 20341
rect 1434 20265 1542 20341
rect 2202 20265 2310 20341
rect 2682 20265 2790 20341
rect 3450 20265 3558 20341
rect 3930 20265 4038 20341
rect 4698 20265 4806 20341
rect 5178 20265 5286 20341
rect 5946 20265 6054 20341
rect 6426 20265 6534 20341
rect 7194 20265 7302 20341
rect 7674 20265 7782 20341
rect 8442 20265 8550 20341
rect 8922 20265 9030 20341
rect 9690 20265 9798 20341
rect 10170 20265 10278 20341
rect 10938 20265 11046 20341
rect 11418 20265 11526 20341
rect 12186 20265 12294 20341
rect 12666 20265 12774 20341
rect 13434 20265 13542 20341
rect 13914 20265 14022 20341
rect 14682 20265 14790 20341
rect 15162 20265 15270 20341
rect 15930 20265 16038 20341
rect 16410 20265 16518 20341
rect 17178 20265 17286 20341
rect 17658 20265 17766 20341
rect 18426 20265 18534 20341
rect 18906 20265 19014 20341
rect 19674 20265 19782 20341
rect 0 20169 19968 20217
rect 0 20073 19968 20121
rect 186 19949 294 20025
rect 954 19949 1062 20025
rect 1434 19949 1542 20025
rect 2202 19949 2310 20025
rect 2682 19949 2790 20025
rect 3450 19949 3558 20025
rect 3930 19949 4038 20025
rect 4698 19949 4806 20025
rect 5178 19949 5286 20025
rect 5946 19949 6054 20025
rect 6426 19949 6534 20025
rect 7194 19949 7302 20025
rect 7674 19949 7782 20025
rect 8442 19949 8550 20025
rect 8922 19949 9030 20025
rect 9690 19949 9798 20025
rect 10170 19949 10278 20025
rect 10938 19949 11046 20025
rect 11418 19949 11526 20025
rect 12186 19949 12294 20025
rect 12666 19949 12774 20025
rect 13434 19949 13542 20025
rect 13914 19949 14022 20025
rect 14682 19949 14790 20025
rect 15162 19949 15270 20025
rect 15930 19949 16038 20025
rect 16410 19949 16518 20025
rect 17178 19949 17286 20025
rect 17658 19949 17766 20025
rect 18426 19949 18534 20025
rect 18906 19949 19014 20025
rect 19674 19949 19782 20025
rect 0 19853 19968 19901
rect 186 19695 294 19805
rect 954 19695 1062 19805
rect 1434 19695 1542 19805
rect 2202 19695 2310 19805
rect 2682 19695 2790 19805
rect 3450 19695 3558 19805
rect 3930 19695 4038 19805
rect 4698 19695 4806 19805
rect 5178 19695 5286 19805
rect 5946 19695 6054 19805
rect 6426 19695 6534 19805
rect 7194 19695 7302 19805
rect 7674 19695 7782 19805
rect 8442 19695 8550 19805
rect 8922 19695 9030 19805
rect 9690 19695 9798 19805
rect 10170 19695 10278 19805
rect 10938 19695 11046 19805
rect 11418 19695 11526 19805
rect 12186 19695 12294 19805
rect 12666 19695 12774 19805
rect 13434 19695 13542 19805
rect 13914 19695 14022 19805
rect 14682 19695 14790 19805
rect 15162 19695 15270 19805
rect 15930 19695 16038 19805
rect 16410 19695 16518 19805
rect 17178 19695 17286 19805
rect 17658 19695 17766 19805
rect 18426 19695 18534 19805
rect 18906 19695 19014 19805
rect 19674 19695 19782 19805
rect 0 19599 19968 19647
rect 186 19475 294 19551
rect 954 19475 1062 19551
rect 1434 19475 1542 19551
rect 2202 19475 2310 19551
rect 2682 19475 2790 19551
rect 3450 19475 3558 19551
rect 3930 19475 4038 19551
rect 4698 19475 4806 19551
rect 5178 19475 5286 19551
rect 5946 19475 6054 19551
rect 6426 19475 6534 19551
rect 7194 19475 7302 19551
rect 7674 19475 7782 19551
rect 8442 19475 8550 19551
rect 8922 19475 9030 19551
rect 9690 19475 9798 19551
rect 10170 19475 10278 19551
rect 10938 19475 11046 19551
rect 11418 19475 11526 19551
rect 12186 19475 12294 19551
rect 12666 19475 12774 19551
rect 13434 19475 13542 19551
rect 13914 19475 14022 19551
rect 14682 19475 14790 19551
rect 15162 19475 15270 19551
rect 15930 19475 16038 19551
rect 16410 19475 16518 19551
rect 17178 19475 17286 19551
rect 17658 19475 17766 19551
rect 18426 19475 18534 19551
rect 18906 19475 19014 19551
rect 19674 19475 19782 19551
rect 0 19379 19968 19427
rect 0 19283 19968 19331
rect 186 19159 294 19235
rect 954 19159 1062 19235
rect 1434 19159 1542 19235
rect 2202 19159 2310 19235
rect 2682 19159 2790 19235
rect 3450 19159 3558 19235
rect 3930 19159 4038 19235
rect 4698 19159 4806 19235
rect 5178 19159 5286 19235
rect 5946 19159 6054 19235
rect 6426 19159 6534 19235
rect 7194 19159 7302 19235
rect 7674 19159 7782 19235
rect 8442 19159 8550 19235
rect 8922 19159 9030 19235
rect 9690 19159 9798 19235
rect 10170 19159 10278 19235
rect 10938 19159 11046 19235
rect 11418 19159 11526 19235
rect 12186 19159 12294 19235
rect 12666 19159 12774 19235
rect 13434 19159 13542 19235
rect 13914 19159 14022 19235
rect 14682 19159 14790 19235
rect 15162 19159 15270 19235
rect 15930 19159 16038 19235
rect 16410 19159 16518 19235
rect 17178 19159 17286 19235
rect 17658 19159 17766 19235
rect 18426 19159 18534 19235
rect 18906 19159 19014 19235
rect 19674 19159 19782 19235
rect 0 19063 19968 19111
rect 186 18905 294 19015
rect 954 18905 1062 19015
rect 1434 18905 1542 19015
rect 2202 18905 2310 19015
rect 2682 18905 2790 19015
rect 3450 18905 3558 19015
rect 3930 18905 4038 19015
rect 4698 18905 4806 19015
rect 5178 18905 5286 19015
rect 5946 18905 6054 19015
rect 6426 18905 6534 19015
rect 7194 18905 7302 19015
rect 7674 18905 7782 19015
rect 8442 18905 8550 19015
rect 8922 18905 9030 19015
rect 9690 18905 9798 19015
rect 10170 18905 10278 19015
rect 10938 18905 11046 19015
rect 11418 18905 11526 19015
rect 12186 18905 12294 19015
rect 12666 18905 12774 19015
rect 13434 18905 13542 19015
rect 13914 18905 14022 19015
rect 14682 18905 14790 19015
rect 15162 18905 15270 19015
rect 15930 18905 16038 19015
rect 16410 18905 16518 19015
rect 17178 18905 17286 19015
rect 17658 18905 17766 19015
rect 18426 18905 18534 19015
rect 18906 18905 19014 19015
rect 19674 18905 19782 19015
rect 0 18809 19968 18857
rect 186 18685 294 18761
rect 954 18685 1062 18761
rect 1434 18685 1542 18761
rect 2202 18685 2310 18761
rect 2682 18685 2790 18761
rect 3450 18685 3558 18761
rect 3930 18685 4038 18761
rect 4698 18685 4806 18761
rect 5178 18685 5286 18761
rect 5946 18685 6054 18761
rect 6426 18685 6534 18761
rect 7194 18685 7302 18761
rect 7674 18685 7782 18761
rect 8442 18685 8550 18761
rect 8922 18685 9030 18761
rect 9690 18685 9798 18761
rect 10170 18685 10278 18761
rect 10938 18685 11046 18761
rect 11418 18685 11526 18761
rect 12186 18685 12294 18761
rect 12666 18685 12774 18761
rect 13434 18685 13542 18761
rect 13914 18685 14022 18761
rect 14682 18685 14790 18761
rect 15162 18685 15270 18761
rect 15930 18685 16038 18761
rect 16410 18685 16518 18761
rect 17178 18685 17286 18761
rect 17658 18685 17766 18761
rect 18426 18685 18534 18761
rect 18906 18685 19014 18761
rect 19674 18685 19782 18761
rect 0 18589 19968 18637
rect 0 18493 19968 18541
rect 186 18369 294 18445
rect 954 18369 1062 18445
rect 1434 18369 1542 18445
rect 2202 18369 2310 18445
rect 2682 18369 2790 18445
rect 3450 18369 3558 18445
rect 3930 18369 4038 18445
rect 4698 18369 4806 18445
rect 5178 18369 5286 18445
rect 5946 18369 6054 18445
rect 6426 18369 6534 18445
rect 7194 18369 7302 18445
rect 7674 18369 7782 18445
rect 8442 18369 8550 18445
rect 8922 18369 9030 18445
rect 9690 18369 9798 18445
rect 10170 18369 10278 18445
rect 10938 18369 11046 18445
rect 11418 18369 11526 18445
rect 12186 18369 12294 18445
rect 12666 18369 12774 18445
rect 13434 18369 13542 18445
rect 13914 18369 14022 18445
rect 14682 18369 14790 18445
rect 15162 18369 15270 18445
rect 15930 18369 16038 18445
rect 16410 18369 16518 18445
rect 17178 18369 17286 18445
rect 17658 18369 17766 18445
rect 18426 18369 18534 18445
rect 18906 18369 19014 18445
rect 19674 18369 19782 18445
rect 0 18273 19968 18321
rect 186 18115 294 18225
rect 954 18115 1062 18225
rect 1434 18115 1542 18225
rect 2202 18115 2310 18225
rect 2682 18115 2790 18225
rect 3450 18115 3558 18225
rect 3930 18115 4038 18225
rect 4698 18115 4806 18225
rect 5178 18115 5286 18225
rect 5946 18115 6054 18225
rect 6426 18115 6534 18225
rect 7194 18115 7302 18225
rect 7674 18115 7782 18225
rect 8442 18115 8550 18225
rect 8922 18115 9030 18225
rect 9690 18115 9798 18225
rect 10170 18115 10278 18225
rect 10938 18115 11046 18225
rect 11418 18115 11526 18225
rect 12186 18115 12294 18225
rect 12666 18115 12774 18225
rect 13434 18115 13542 18225
rect 13914 18115 14022 18225
rect 14682 18115 14790 18225
rect 15162 18115 15270 18225
rect 15930 18115 16038 18225
rect 16410 18115 16518 18225
rect 17178 18115 17286 18225
rect 17658 18115 17766 18225
rect 18426 18115 18534 18225
rect 18906 18115 19014 18225
rect 19674 18115 19782 18225
rect 0 18019 19968 18067
rect 186 17895 294 17971
rect 954 17895 1062 17971
rect 1434 17895 1542 17971
rect 2202 17895 2310 17971
rect 2682 17895 2790 17971
rect 3450 17895 3558 17971
rect 3930 17895 4038 17971
rect 4698 17895 4806 17971
rect 5178 17895 5286 17971
rect 5946 17895 6054 17971
rect 6426 17895 6534 17971
rect 7194 17895 7302 17971
rect 7674 17895 7782 17971
rect 8442 17895 8550 17971
rect 8922 17895 9030 17971
rect 9690 17895 9798 17971
rect 10170 17895 10278 17971
rect 10938 17895 11046 17971
rect 11418 17895 11526 17971
rect 12186 17895 12294 17971
rect 12666 17895 12774 17971
rect 13434 17895 13542 17971
rect 13914 17895 14022 17971
rect 14682 17895 14790 17971
rect 15162 17895 15270 17971
rect 15930 17895 16038 17971
rect 16410 17895 16518 17971
rect 17178 17895 17286 17971
rect 17658 17895 17766 17971
rect 18426 17895 18534 17971
rect 18906 17895 19014 17971
rect 19674 17895 19782 17971
rect 0 17799 19968 17847
rect 0 17703 19968 17751
rect 186 17579 294 17655
rect 954 17579 1062 17655
rect 1434 17579 1542 17655
rect 2202 17579 2310 17655
rect 2682 17579 2790 17655
rect 3450 17579 3558 17655
rect 3930 17579 4038 17655
rect 4698 17579 4806 17655
rect 5178 17579 5286 17655
rect 5946 17579 6054 17655
rect 6426 17579 6534 17655
rect 7194 17579 7302 17655
rect 7674 17579 7782 17655
rect 8442 17579 8550 17655
rect 8922 17579 9030 17655
rect 9690 17579 9798 17655
rect 10170 17579 10278 17655
rect 10938 17579 11046 17655
rect 11418 17579 11526 17655
rect 12186 17579 12294 17655
rect 12666 17579 12774 17655
rect 13434 17579 13542 17655
rect 13914 17579 14022 17655
rect 14682 17579 14790 17655
rect 15162 17579 15270 17655
rect 15930 17579 16038 17655
rect 16410 17579 16518 17655
rect 17178 17579 17286 17655
rect 17658 17579 17766 17655
rect 18426 17579 18534 17655
rect 18906 17579 19014 17655
rect 19674 17579 19782 17655
rect 0 17483 19968 17531
rect 186 17325 294 17435
rect 954 17325 1062 17435
rect 1434 17325 1542 17435
rect 2202 17325 2310 17435
rect 2682 17325 2790 17435
rect 3450 17325 3558 17435
rect 3930 17325 4038 17435
rect 4698 17325 4806 17435
rect 5178 17325 5286 17435
rect 5946 17325 6054 17435
rect 6426 17325 6534 17435
rect 7194 17325 7302 17435
rect 7674 17325 7782 17435
rect 8442 17325 8550 17435
rect 8922 17325 9030 17435
rect 9690 17325 9798 17435
rect 10170 17325 10278 17435
rect 10938 17325 11046 17435
rect 11418 17325 11526 17435
rect 12186 17325 12294 17435
rect 12666 17325 12774 17435
rect 13434 17325 13542 17435
rect 13914 17325 14022 17435
rect 14682 17325 14790 17435
rect 15162 17325 15270 17435
rect 15930 17325 16038 17435
rect 16410 17325 16518 17435
rect 17178 17325 17286 17435
rect 17658 17325 17766 17435
rect 18426 17325 18534 17435
rect 18906 17325 19014 17435
rect 19674 17325 19782 17435
rect 0 17229 19968 17277
rect 186 17105 294 17181
rect 954 17105 1062 17181
rect 1434 17105 1542 17181
rect 2202 17105 2310 17181
rect 2682 17105 2790 17181
rect 3450 17105 3558 17181
rect 3930 17105 4038 17181
rect 4698 17105 4806 17181
rect 5178 17105 5286 17181
rect 5946 17105 6054 17181
rect 6426 17105 6534 17181
rect 7194 17105 7302 17181
rect 7674 17105 7782 17181
rect 8442 17105 8550 17181
rect 8922 17105 9030 17181
rect 9690 17105 9798 17181
rect 10170 17105 10278 17181
rect 10938 17105 11046 17181
rect 11418 17105 11526 17181
rect 12186 17105 12294 17181
rect 12666 17105 12774 17181
rect 13434 17105 13542 17181
rect 13914 17105 14022 17181
rect 14682 17105 14790 17181
rect 15162 17105 15270 17181
rect 15930 17105 16038 17181
rect 16410 17105 16518 17181
rect 17178 17105 17286 17181
rect 17658 17105 17766 17181
rect 18426 17105 18534 17181
rect 18906 17105 19014 17181
rect 19674 17105 19782 17181
rect 0 17009 19968 17057
rect 0 16913 19968 16961
rect 186 16789 294 16865
rect 954 16789 1062 16865
rect 1434 16789 1542 16865
rect 2202 16789 2310 16865
rect 2682 16789 2790 16865
rect 3450 16789 3558 16865
rect 3930 16789 4038 16865
rect 4698 16789 4806 16865
rect 5178 16789 5286 16865
rect 5946 16789 6054 16865
rect 6426 16789 6534 16865
rect 7194 16789 7302 16865
rect 7674 16789 7782 16865
rect 8442 16789 8550 16865
rect 8922 16789 9030 16865
rect 9690 16789 9798 16865
rect 10170 16789 10278 16865
rect 10938 16789 11046 16865
rect 11418 16789 11526 16865
rect 12186 16789 12294 16865
rect 12666 16789 12774 16865
rect 13434 16789 13542 16865
rect 13914 16789 14022 16865
rect 14682 16789 14790 16865
rect 15162 16789 15270 16865
rect 15930 16789 16038 16865
rect 16410 16789 16518 16865
rect 17178 16789 17286 16865
rect 17658 16789 17766 16865
rect 18426 16789 18534 16865
rect 18906 16789 19014 16865
rect 19674 16789 19782 16865
rect 0 16693 19968 16741
rect 186 16535 294 16645
rect 954 16535 1062 16645
rect 1434 16535 1542 16645
rect 2202 16535 2310 16645
rect 2682 16535 2790 16645
rect 3450 16535 3558 16645
rect 3930 16535 4038 16645
rect 4698 16535 4806 16645
rect 5178 16535 5286 16645
rect 5946 16535 6054 16645
rect 6426 16535 6534 16645
rect 7194 16535 7302 16645
rect 7674 16535 7782 16645
rect 8442 16535 8550 16645
rect 8922 16535 9030 16645
rect 9690 16535 9798 16645
rect 10170 16535 10278 16645
rect 10938 16535 11046 16645
rect 11418 16535 11526 16645
rect 12186 16535 12294 16645
rect 12666 16535 12774 16645
rect 13434 16535 13542 16645
rect 13914 16535 14022 16645
rect 14682 16535 14790 16645
rect 15162 16535 15270 16645
rect 15930 16535 16038 16645
rect 16410 16535 16518 16645
rect 17178 16535 17286 16645
rect 17658 16535 17766 16645
rect 18426 16535 18534 16645
rect 18906 16535 19014 16645
rect 19674 16535 19782 16645
rect 0 16439 19968 16487
rect 186 16315 294 16391
rect 954 16315 1062 16391
rect 1434 16315 1542 16391
rect 2202 16315 2310 16391
rect 2682 16315 2790 16391
rect 3450 16315 3558 16391
rect 3930 16315 4038 16391
rect 4698 16315 4806 16391
rect 5178 16315 5286 16391
rect 5946 16315 6054 16391
rect 6426 16315 6534 16391
rect 7194 16315 7302 16391
rect 7674 16315 7782 16391
rect 8442 16315 8550 16391
rect 8922 16315 9030 16391
rect 9690 16315 9798 16391
rect 10170 16315 10278 16391
rect 10938 16315 11046 16391
rect 11418 16315 11526 16391
rect 12186 16315 12294 16391
rect 12666 16315 12774 16391
rect 13434 16315 13542 16391
rect 13914 16315 14022 16391
rect 14682 16315 14790 16391
rect 15162 16315 15270 16391
rect 15930 16315 16038 16391
rect 16410 16315 16518 16391
rect 17178 16315 17286 16391
rect 17658 16315 17766 16391
rect 18426 16315 18534 16391
rect 18906 16315 19014 16391
rect 19674 16315 19782 16391
rect 0 16219 19968 16267
rect 0 16123 19968 16171
rect 186 15999 294 16075
rect 954 15999 1062 16075
rect 1434 15999 1542 16075
rect 2202 15999 2310 16075
rect 2682 15999 2790 16075
rect 3450 15999 3558 16075
rect 3930 15999 4038 16075
rect 4698 15999 4806 16075
rect 5178 15999 5286 16075
rect 5946 15999 6054 16075
rect 6426 15999 6534 16075
rect 7194 15999 7302 16075
rect 7674 15999 7782 16075
rect 8442 15999 8550 16075
rect 8922 15999 9030 16075
rect 9690 15999 9798 16075
rect 10170 15999 10278 16075
rect 10938 15999 11046 16075
rect 11418 15999 11526 16075
rect 12186 15999 12294 16075
rect 12666 15999 12774 16075
rect 13434 15999 13542 16075
rect 13914 15999 14022 16075
rect 14682 15999 14790 16075
rect 15162 15999 15270 16075
rect 15930 15999 16038 16075
rect 16410 15999 16518 16075
rect 17178 15999 17286 16075
rect 17658 15999 17766 16075
rect 18426 15999 18534 16075
rect 18906 15999 19014 16075
rect 19674 15999 19782 16075
rect 0 15903 19968 15951
rect 186 15745 294 15855
rect 954 15745 1062 15855
rect 1434 15745 1542 15855
rect 2202 15745 2310 15855
rect 2682 15745 2790 15855
rect 3450 15745 3558 15855
rect 3930 15745 4038 15855
rect 4698 15745 4806 15855
rect 5178 15745 5286 15855
rect 5946 15745 6054 15855
rect 6426 15745 6534 15855
rect 7194 15745 7302 15855
rect 7674 15745 7782 15855
rect 8442 15745 8550 15855
rect 8922 15745 9030 15855
rect 9690 15745 9798 15855
rect 10170 15745 10278 15855
rect 10938 15745 11046 15855
rect 11418 15745 11526 15855
rect 12186 15745 12294 15855
rect 12666 15745 12774 15855
rect 13434 15745 13542 15855
rect 13914 15745 14022 15855
rect 14682 15745 14790 15855
rect 15162 15745 15270 15855
rect 15930 15745 16038 15855
rect 16410 15745 16518 15855
rect 17178 15745 17286 15855
rect 17658 15745 17766 15855
rect 18426 15745 18534 15855
rect 18906 15745 19014 15855
rect 19674 15745 19782 15855
rect 0 15649 19968 15697
rect 186 15525 294 15601
rect 954 15525 1062 15601
rect 1434 15525 1542 15601
rect 2202 15525 2310 15601
rect 2682 15525 2790 15601
rect 3450 15525 3558 15601
rect 3930 15525 4038 15601
rect 4698 15525 4806 15601
rect 5178 15525 5286 15601
rect 5946 15525 6054 15601
rect 6426 15525 6534 15601
rect 7194 15525 7302 15601
rect 7674 15525 7782 15601
rect 8442 15525 8550 15601
rect 8922 15525 9030 15601
rect 9690 15525 9798 15601
rect 10170 15525 10278 15601
rect 10938 15525 11046 15601
rect 11418 15525 11526 15601
rect 12186 15525 12294 15601
rect 12666 15525 12774 15601
rect 13434 15525 13542 15601
rect 13914 15525 14022 15601
rect 14682 15525 14790 15601
rect 15162 15525 15270 15601
rect 15930 15525 16038 15601
rect 16410 15525 16518 15601
rect 17178 15525 17286 15601
rect 17658 15525 17766 15601
rect 18426 15525 18534 15601
rect 18906 15525 19014 15601
rect 19674 15525 19782 15601
rect 0 15429 19968 15477
rect 0 15333 19968 15381
rect 186 15209 294 15285
rect 954 15209 1062 15285
rect 1434 15209 1542 15285
rect 2202 15209 2310 15285
rect 2682 15209 2790 15285
rect 3450 15209 3558 15285
rect 3930 15209 4038 15285
rect 4698 15209 4806 15285
rect 5178 15209 5286 15285
rect 5946 15209 6054 15285
rect 6426 15209 6534 15285
rect 7194 15209 7302 15285
rect 7674 15209 7782 15285
rect 8442 15209 8550 15285
rect 8922 15209 9030 15285
rect 9690 15209 9798 15285
rect 10170 15209 10278 15285
rect 10938 15209 11046 15285
rect 11418 15209 11526 15285
rect 12186 15209 12294 15285
rect 12666 15209 12774 15285
rect 13434 15209 13542 15285
rect 13914 15209 14022 15285
rect 14682 15209 14790 15285
rect 15162 15209 15270 15285
rect 15930 15209 16038 15285
rect 16410 15209 16518 15285
rect 17178 15209 17286 15285
rect 17658 15209 17766 15285
rect 18426 15209 18534 15285
rect 18906 15209 19014 15285
rect 19674 15209 19782 15285
rect 0 15113 19968 15161
rect 186 14955 294 15065
rect 954 14955 1062 15065
rect 1434 14955 1542 15065
rect 2202 14955 2310 15065
rect 2682 14955 2790 15065
rect 3450 14955 3558 15065
rect 3930 14955 4038 15065
rect 4698 14955 4806 15065
rect 5178 14955 5286 15065
rect 5946 14955 6054 15065
rect 6426 14955 6534 15065
rect 7194 14955 7302 15065
rect 7674 14955 7782 15065
rect 8442 14955 8550 15065
rect 8922 14955 9030 15065
rect 9690 14955 9798 15065
rect 10170 14955 10278 15065
rect 10938 14955 11046 15065
rect 11418 14955 11526 15065
rect 12186 14955 12294 15065
rect 12666 14955 12774 15065
rect 13434 14955 13542 15065
rect 13914 14955 14022 15065
rect 14682 14955 14790 15065
rect 15162 14955 15270 15065
rect 15930 14955 16038 15065
rect 16410 14955 16518 15065
rect 17178 14955 17286 15065
rect 17658 14955 17766 15065
rect 18426 14955 18534 15065
rect 18906 14955 19014 15065
rect 19674 14955 19782 15065
rect 0 14859 19968 14907
rect 186 14735 294 14811
rect 954 14735 1062 14811
rect 1434 14735 1542 14811
rect 2202 14735 2310 14811
rect 2682 14735 2790 14811
rect 3450 14735 3558 14811
rect 3930 14735 4038 14811
rect 4698 14735 4806 14811
rect 5178 14735 5286 14811
rect 5946 14735 6054 14811
rect 6426 14735 6534 14811
rect 7194 14735 7302 14811
rect 7674 14735 7782 14811
rect 8442 14735 8550 14811
rect 8922 14735 9030 14811
rect 9690 14735 9798 14811
rect 10170 14735 10278 14811
rect 10938 14735 11046 14811
rect 11418 14735 11526 14811
rect 12186 14735 12294 14811
rect 12666 14735 12774 14811
rect 13434 14735 13542 14811
rect 13914 14735 14022 14811
rect 14682 14735 14790 14811
rect 15162 14735 15270 14811
rect 15930 14735 16038 14811
rect 16410 14735 16518 14811
rect 17178 14735 17286 14811
rect 17658 14735 17766 14811
rect 18426 14735 18534 14811
rect 18906 14735 19014 14811
rect 19674 14735 19782 14811
rect 0 14639 19968 14687
rect 0 14543 19968 14591
rect 186 14419 294 14495
rect 954 14419 1062 14495
rect 1434 14419 1542 14495
rect 2202 14419 2310 14495
rect 2682 14419 2790 14495
rect 3450 14419 3558 14495
rect 3930 14419 4038 14495
rect 4698 14419 4806 14495
rect 5178 14419 5286 14495
rect 5946 14419 6054 14495
rect 6426 14419 6534 14495
rect 7194 14419 7302 14495
rect 7674 14419 7782 14495
rect 8442 14419 8550 14495
rect 8922 14419 9030 14495
rect 9690 14419 9798 14495
rect 10170 14419 10278 14495
rect 10938 14419 11046 14495
rect 11418 14419 11526 14495
rect 12186 14419 12294 14495
rect 12666 14419 12774 14495
rect 13434 14419 13542 14495
rect 13914 14419 14022 14495
rect 14682 14419 14790 14495
rect 15162 14419 15270 14495
rect 15930 14419 16038 14495
rect 16410 14419 16518 14495
rect 17178 14419 17286 14495
rect 17658 14419 17766 14495
rect 18426 14419 18534 14495
rect 18906 14419 19014 14495
rect 19674 14419 19782 14495
rect 0 14323 19968 14371
rect 186 14165 294 14275
rect 954 14165 1062 14275
rect 1434 14165 1542 14275
rect 2202 14165 2310 14275
rect 2682 14165 2790 14275
rect 3450 14165 3558 14275
rect 3930 14165 4038 14275
rect 4698 14165 4806 14275
rect 5178 14165 5286 14275
rect 5946 14165 6054 14275
rect 6426 14165 6534 14275
rect 7194 14165 7302 14275
rect 7674 14165 7782 14275
rect 8442 14165 8550 14275
rect 8922 14165 9030 14275
rect 9690 14165 9798 14275
rect 10170 14165 10278 14275
rect 10938 14165 11046 14275
rect 11418 14165 11526 14275
rect 12186 14165 12294 14275
rect 12666 14165 12774 14275
rect 13434 14165 13542 14275
rect 13914 14165 14022 14275
rect 14682 14165 14790 14275
rect 15162 14165 15270 14275
rect 15930 14165 16038 14275
rect 16410 14165 16518 14275
rect 17178 14165 17286 14275
rect 17658 14165 17766 14275
rect 18426 14165 18534 14275
rect 18906 14165 19014 14275
rect 19674 14165 19782 14275
rect 0 14069 19968 14117
rect 186 13945 294 14021
rect 954 13945 1062 14021
rect 1434 13945 1542 14021
rect 2202 13945 2310 14021
rect 2682 13945 2790 14021
rect 3450 13945 3558 14021
rect 3930 13945 4038 14021
rect 4698 13945 4806 14021
rect 5178 13945 5286 14021
rect 5946 13945 6054 14021
rect 6426 13945 6534 14021
rect 7194 13945 7302 14021
rect 7674 13945 7782 14021
rect 8442 13945 8550 14021
rect 8922 13945 9030 14021
rect 9690 13945 9798 14021
rect 10170 13945 10278 14021
rect 10938 13945 11046 14021
rect 11418 13945 11526 14021
rect 12186 13945 12294 14021
rect 12666 13945 12774 14021
rect 13434 13945 13542 14021
rect 13914 13945 14022 14021
rect 14682 13945 14790 14021
rect 15162 13945 15270 14021
rect 15930 13945 16038 14021
rect 16410 13945 16518 14021
rect 17178 13945 17286 14021
rect 17658 13945 17766 14021
rect 18426 13945 18534 14021
rect 18906 13945 19014 14021
rect 19674 13945 19782 14021
rect 0 13849 19968 13897
rect 0 13753 19968 13801
rect 186 13629 294 13705
rect 954 13629 1062 13705
rect 1434 13629 1542 13705
rect 2202 13629 2310 13705
rect 2682 13629 2790 13705
rect 3450 13629 3558 13705
rect 3930 13629 4038 13705
rect 4698 13629 4806 13705
rect 5178 13629 5286 13705
rect 5946 13629 6054 13705
rect 6426 13629 6534 13705
rect 7194 13629 7302 13705
rect 7674 13629 7782 13705
rect 8442 13629 8550 13705
rect 8922 13629 9030 13705
rect 9690 13629 9798 13705
rect 10170 13629 10278 13705
rect 10938 13629 11046 13705
rect 11418 13629 11526 13705
rect 12186 13629 12294 13705
rect 12666 13629 12774 13705
rect 13434 13629 13542 13705
rect 13914 13629 14022 13705
rect 14682 13629 14790 13705
rect 15162 13629 15270 13705
rect 15930 13629 16038 13705
rect 16410 13629 16518 13705
rect 17178 13629 17286 13705
rect 17658 13629 17766 13705
rect 18426 13629 18534 13705
rect 18906 13629 19014 13705
rect 19674 13629 19782 13705
rect 0 13533 19968 13581
rect 186 13375 294 13485
rect 954 13375 1062 13485
rect 1434 13375 1542 13485
rect 2202 13375 2310 13485
rect 2682 13375 2790 13485
rect 3450 13375 3558 13485
rect 3930 13375 4038 13485
rect 4698 13375 4806 13485
rect 5178 13375 5286 13485
rect 5946 13375 6054 13485
rect 6426 13375 6534 13485
rect 7194 13375 7302 13485
rect 7674 13375 7782 13485
rect 8442 13375 8550 13485
rect 8922 13375 9030 13485
rect 9690 13375 9798 13485
rect 10170 13375 10278 13485
rect 10938 13375 11046 13485
rect 11418 13375 11526 13485
rect 12186 13375 12294 13485
rect 12666 13375 12774 13485
rect 13434 13375 13542 13485
rect 13914 13375 14022 13485
rect 14682 13375 14790 13485
rect 15162 13375 15270 13485
rect 15930 13375 16038 13485
rect 16410 13375 16518 13485
rect 17178 13375 17286 13485
rect 17658 13375 17766 13485
rect 18426 13375 18534 13485
rect 18906 13375 19014 13485
rect 19674 13375 19782 13485
rect 0 13279 19968 13327
rect 186 13155 294 13231
rect 954 13155 1062 13231
rect 1434 13155 1542 13231
rect 2202 13155 2310 13231
rect 2682 13155 2790 13231
rect 3450 13155 3558 13231
rect 3930 13155 4038 13231
rect 4698 13155 4806 13231
rect 5178 13155 5286 13231
rect 5946 13155 6054 13231
rect 6426 13155 6534 13231
rect 7194 13155 7302 13231
rect 7674 13155 7782 13231
rect 8442 13155 8550 13231
rect 8922 13155 9030 13231
rect 9690 13155 9798 13231
rect 10170 13155 10278 13231
rect 10938 13155 11046 13231
rect 11418 13155 11526 13231
rect 12186 13155 12294 13231
rect 12666 13155 12774 13231
rect 13434 13155 13542 13231
rect 13914 13155 14022 13231
rect 14682 13155 14790 13231
rect 15162 13155 15270 13231
rect 15930 13155 16038 13231
rect 16410 13155 16518 13231
rect 17178 13155 17286 13231
rect 17658 13155 17766 13231
rect 18426 13155 18534 13231
rect 18906 13155 19014 13231
rect 19674 13155 19782 13231
rect 0 13059 19968 13107
rect 0 12963 19968 13011
rect 186 12839 294 12915
rect 954 12839 1062 12915
rect 1434 12839 1542 12915
rect 2202 12839 2310 12915
rect 2682 12839 2790 12915
rect 3450 12839 3558 12915
rect 3930 12839 4038 12915
rect 4698 12839 4806 12915
rect 5178 12839 5286 12915
rect 5946 12839 6054 12915
rect 6426 12839 6534 12915
rect 7194 12839 7302 12915
rect 7674 12839 7782 12915
rect 8442 12839 8550 12915
rect 8922 12839 9030 12915
rect 9690 12839 9798 12915
rect 10170 12839 10278 12915
rect 10938 12839 11046 12915
rect 11418 12839 11526 12915
rect 12186 12839 12294 12915
rect 12666 12839 12774 12915
rect 13434 12839 13542 12915
rect 13914 12839 14022 12915
rect 14682 12839 14790 12915
rect 15162 12839 15270 12915
rect 15930 12839 16038 12915
rect 16410 12839 16518 12915
rect 17178 12839 17286 12915
rect 17658 12839 17766 12915
rect 18426 12839 18534 12915
rect 18906 12839 19014 12915
rect 19674 12839 19782 12915
rect 0 12743 19968 12791
rect 186 12585 294 12695
rect 954 12585 1062 12695
rect 1434 12585 1542 12695
rect 2202 12585 2310 12695
rect 2682 12585 2790 12695
rect 3450 12585 3558 12695
rect 3930 12585 4038 12695
rect 4698 12585 4806 12695
rect 5178 12585 5286 12695
rect 5946 12585 6054 12695
rect 6426 12585 6534 12695
rect 7194 12585 7302 12695
rect 7674 12585 7782 12695
rect 8442 12585 8550 12695
rect 8922 12585 9030 12695
rect 9690 12585 9798 12695
rect 10170 12585 10278 12695
rect 10938 12585 11046 12695
rect 11418 12585 11526 12695
rect 12186 12585 12294 12695
rect 12666 12585 12774 12695
rect 13434 12585 13542 12695
rect 13914 12585 14022 12695
rect 14682 12585 14790 12695
rect 15162 12585 15270 12695
rect 15930 12585 16038 12695
rect 16410 12585 16518 12695
rect 17178 12585 17286 12695
rect 17658 12585 17766 12695
rect 18426 12585 18534 12695
rect 18906 12585 19014 12695
rect 19674 12585 19782 12695
rect 0 12489 19968 12537
rect 186 12365 294 12441
rect 954 12365 1062 12441
rect 1434 12365 1542 12441
rect 2202 12365 2310 12441
rect 2682 12365 2790 12441
rect 3450 12365 3558 12441
rect 3930 12365 4038 12441
rect 4698 12365 4806 12441
rect 5178 12365 5286 12441
rect 5946 12365 6054 12441
rect 6426 12365 6534 12441
rect 7194 12365 7302 12441
rect 7674 12365 7782 12441
rect 8442 12365 8550 12441
rect 8922 12365 9030 12441
rect 9690 12365 9798 12441
rect 10170 12365 10278 12441
rect 10938 12365 11046 12441
rect 11418 12365 11526 12441
rect 12186 12365 12294 12441
rect 12666 12365 12774 12441
rect 13434 12365 13542 12441
rect 13914 12365 14022 12441
rect 14682 12365 14790 12441
rect 15162 12365 15270 12441
rect 15930 12365 16038 12441
rect 16410 12365 16518 12441
rect 17178 12365 17286 12441
rect 17658 12365 17766 12441
rect 18426 12365 18534 12441
rect 18906 12365 19014 12441
rect 19674 12365 19782 12441
rect 0 12269 19968 12317
rect 0 12173 19968 12221
rect 186 12049 294 12125
rect 954 12049 1062 12125
rect 1434 12049 1542 12125
rect 2202 12049 2310 12125
rect 2682 12049 2790 12125
rect 3450 12049 3558 12125
rect 3930 12049 4038 12125
rect 4698 12049 4806 12125
rect 5178 12049 5286 12125
rect 5946 12049 6054 12125
rect 6426 12049 6534 12125
rect 7194 12049 7302 12125
rect 7674 12049 7782 12125
rect 8442 12049 8550 12125
rect 8922 12049 9030 12125
rect 9690 12049 9798 12125
rect 10170 12049 10278 12125
rect 10938 12049 11046 12125
rect 11418 12049 11526 12125
rect 12186 12049 12294 12125
rect 12666 12049 12774 12125
rect 13434 12049 13542 12125
rect 13914 12049 14022 12125
rect 14682 12049 14790 12125
rect 15162 12049 15270 12125
rect 15930 12049 16038 12125
rect 16410 12049 16518 12125
rect 17178 12049 17286 12125
rect 17658 12049 17766 12125
rect 18426 12049 18534 12125
rect 18906 12049 19014 12125
rect 19674 12049 19782 12125
rect 0 11953 19968 12001
rect 186 11795 294 11905
rect 954 11795 1062 11905
rect 1434 11795 1542 11905
rect 2202 11795 2310 11905
rect 2682 11795 2790 11905
rect 3450 11795 3558 11905
rect 3930 11795 4038 11905
rect 4698 11795 4806 11905
rect 5178 11795 5286 11905
rect 5946 11795 6054 11905
rect 6426 11795 6534 11905
rect 7194 11795 7302 11905
rect 7674 11795 7782 11905
rect 8442 11795 8550 11905
rect 8922 11795 9030 11905
rect 9690 11795 9798 11905
rect 10170 11795 10278 11905
rect 10938 11795 11046 11905
rect 11418 11795 11526 11905
rect 12186 11795 12294 11905
rect 12666 11795 12774 11905
rect 13434 11795 13542 11905
rect 13914 11795 14022 11905
rect 14682 11795 14790 11905
rect 15162 11795 15270 11905
rect 15930 11795 16038 11905
rect 16410 11795 16518 11905
rect 17178 11795 17286 11905
rect 17658 11795 17766 11905
rect 18426 11795 18534 11905
rect 18906 11795 19014 11905
rect 19674 11795 19782 11905
rect 0 11699 19968 11747
rect 186 11575 294 11651
rect 954 11575 1062 11651
rect 1434 11575 1542 11651
rect 2202 11575 2310 11651
rect 2682 11575 2790 11651
rect 3450 11575 3558 11651
rect 3930 11575 4038 11651
rect 4698 11575 4806 11651
rect 5178 11575 5286 11651
rect 5946 11575 6054 11651
rect 6426 11575 6534 11651
rect 7194 11575 7302 11651
rect 7674 11575 7782 11651
rect 8442 11575 8550 11651
rect 8922 11575 9030 11651
rect 9690 11575 9798 11651
rect 10170 11575 10278 11651
rect 10938 11575 11046 11651
rect 11418 11575 11526 11651
rect 12186 11575 12294 11651
rect 12666 11575 12774 11651
rect 13434 11575 13542 11651
rect 13914 11575 14022 11651
rect 14682 11575 14790 11651
rect 15162 11575 15270 11651
rect 15930 11575 16038 11651
rect 16410 11575 16518 11651
rect 17178 11575 17286 11651
rect 17658 11575 17766 11651
rect 18426 11575 18534 11651
rect 18906 11575 19014 11651
rect 19674 11575 19782 11651
rect 0 11479 19968 11527
rect 0 11383 19968 11431
rect 186 11259 294 11335
rect 954 11259 1062 11335
rect 1434 11259 1542 11335
rect 2202 11259 2310 11335
rect 2682 11259 2790 11335
rect 3450 11259 3558 11335
rect 3930 11259 4038 11335
rect 4698 11259 4806 11335
rect 5178 11259 5286 11335
rect 5946 11259 6054 11335
rect 6426 11259 6534 11335
rect 7194 11259 7302 11335
rect 7674 11259 7782 11335
rect 8442 11259 8550 11335
rect 8922 11259 9030 11335
rect 9690 11259 9798 11335
rect 10170 11259 10278 11335
rect 10938 11259 11046 11335
rect 11418 11259 11526 11335
rect 12186 11259 12294 11335
rect 12666 11259 12774 11335
rect 13434 11259 13542 11335
rect 13914 11259 14022 11335
rect 14682 11259 14790 11335
rect 15162 11259 15270 11335
rect 15930 11259 16038 11335
rect 16410 11259 16518 11335
rect 17178 11259 17286 11335
rect 17658 11259 17766 11335
rect 18426 11259 18534 11335
rect 18906 11259 19014 11335
rect 19674 11259 19782 11335
rect 0 11163 19968 11211
rect 186 11005 294 11115
rect 954 11005 1062 11115
rect 1434 11005 1542 11115
rect 2202 11005 2310 11115
rect 2682 11005 2790 11115
rect 3450 11005 3558 11115
rect 3930 11005 4038 11115
rect 4698 11005 4806 11115
rect 5178 11005 5286 11115
rect 5946 11005 6054 11115
rect 6426 11005 6534 11115
rect 7194 11005 7302 11115
rect 7674 11005 7782 11115
rect 8442 11005 8550 11115
rect 8922 11005 9030 11115
rect 9690 11005 9798 11115
rect 10170 11005 10278 11115
rect 10938 11005 11046 11115
rect 11418 11005 11526 11115
rect 12186 11005 12294 11115
rect 12666 11005 12774 11115
rect 13434 11005 13542 11115
rect 13914 11005 14022 11115
rect 14682 11005 14790 11115
rect 15162 11005 15270 11115
rect 15930 11005 16038 11115
rect 16410 11005 16518 11115
rect 17178 11005 17286 11115
rect 17658 11005 17766 11115
rect 18426 11005 18534 11115
rect 18906 11005 19014 11115
rect 19674 11005 19782 11115
rect 0 10909 19968 10957
rect 186 10785 294 10861
rect 954 10785 1062 10861
rect 1434 10785 1542 10861
rect 2202 10785 2310 10861
rect 2682 10785 2790 10861
rect 3450 10785 3558 10861
rect 3930 10785 4038 10861
rect 4698 10785 4806 10861
rect 5178 10785 5286 10861
rect 5946 10785 6054 10861
rect 6426 10785 6534 10861
rect 7194 10785 7302 10861
rect 7674 10785 7782 10861
rect 8442 10785 8550 10861
rect 8922 10785 9030 10861
rect 9690 10785 9798 10861
rect 10170 10785 10278 10861
rect 10938 10785 11046 10861
rect 11418 10785 11526 10861
rect 12186 10785 12294 10861
rect 12666 10785 12774 10861
rect 13434 10785 13542 10861
rect 13914 10785 14022 10861
rect 14682 10785 14790 10861
rect 15162 10785 15270 10861
rect 15930 10785 16038 10861
rect 16410 10785 16518 10861
rect 17178 10785 17286 10861
rect 17658 10785 17766 10861
rect 18426 10785 18534 10861
rect 18906 10785 19014 10861
rect 19674 10785 19782 10861
rect 0 10689 19968 10737
rect 0 10593 19968 10641
rect 186 10469 294 10545
rect 954 10469 1062 10545
rect 1434 10469 1542 10545
rect 2202 10469 2310 10545
rect 2682 10469 2790 10545
rect 3450 10469 3558 10545
rect 3930 10469 4038 10545
rect 4698 10469 4806 10545
rect 5178 10469 5286 10545
rect 5946 10469 6054 10545
rect 6426 10469 6534 10545
rect 7194 10469 7302 10545
rect 7674 10469 7782 10545
rect 8442 10469 8550 10545
rect 8922 10469 9030 10545
rect 9690 10469 9798 10545
rect 10170 10469 10278 10545
rect 10938 10469 11046 10545
rect 11418 10469 11526 10545
rect 12186 10469 12294 10545
rect 12666 10469 12774 10545
rect 13434 10469 13542 10545
rect 13914 10469 14022 10545
rect 14682 10469 14790 10545
rect 15162 10469 15270 10545
rect 15930 10469 16038 10545
rect 16410 10469 16518 10545
rect 17178 10469 17286 10545
rect 17658 10469 17766 10545
rect 18426 10469 18534 10545
rect 18906 10469 19014 10545
rect 19674 10469 19782 10545
rect 0 10373 19968 10421
rect 186 10215 294 10325
rect 954 10215 1062 10325
rect 1434 10215 1542 10325
rect 2202 10215 2310 10325
rect 2682 10215 2790 10325
rect 3450 10215 3558 10325
rect 3930 10215 4038 10325
rect 4698 10215 4806 10325
rect 5178 10215 5286 10325
rect 5946 10215 6054 10325
rect 6426 10215 6534 10325
rect 7194 10215 7302 10325
rect 7674 10215 7782 10325
rect 8442 10215 8550 10325
rect 8922 10215 9030 10325
rect 9690 10215 9798 10325
rect 10170 10215 10278 10325
rect 10938 10215 11046 10325
rect 11418 10215 11526 10325
rect 12186 10215 12294 10325
rect 12666 10215 12774 10325
rect 13434 10215 13542 10325
rect 13914 10215 14022 10325
rect 14682 10215 14790 10325
rect 15162 10215 15270 10325
rect 15930 10215 16038 10325
rect 16410 10215 16518 10325
rect 17178 10215 17286 10325
rect 17658 10215 17766 10325
rect 18426 10215 18534 10325
rect 18906 10215 19014 10325
rect 19674 10215 19782 10325
rect 0 10119 19968 10167
rect 186 9995 294 10071
rect 954 9995 1062 10071
rect 1434 9995 1542 10071
rect 2202 9995 2310 10071
rect 2682 9995 2790 10071
rect 3450 9995 3558 10071
rect 3930 9995 4038 10071
rect 4698 9995 4806 10071
rect 5178 9995 5286 10071
rect 5946 9995 6054 10071
rect 6426 9995 6534 10071
rect 7194 9995 7302 10071
rect 7674 9995 7782 10071
rect 8442 9995 8550 10071
rect 8922 9995 9030 10071
rect 9690 9995 9798 10071
rect 10170 9995 10278 10071
rect 10938 9995 11046 10071
rect 11418 9995 11526 10071
rect 12186 9995 12294 10071
rect 12666 9995 12774 10071
rect 13434 9995 13542 10071
rect 13914 9995 14022 10071
rect 14682 9995 14790 10071
rect 15162 9995 15270 10071
rect 15930 9995 16038 10071
rect 16410 9995 16518 10071
rect 17178 9995 17286 10071
rect 17658 9995 17766 10071
rect 18426 9995 18534 10071
rect 18906 9995 19014 10071
rect 19674 9995 19782 10071
rect 0 9899 19968 9947
rect 0 9803 19968 9851
rect 186 9679 294 9755
rect 954 9679 1062 9755
rect 1434 9679 1542 9755
rect 2202 9679 2310 9755
rect 2682 9679 2790 9755
rect 3450 9679 3558 9755
rect 3930 9679 4038 9755
rect 4698 9679 4806 9755
rect 5178 9679 5286 9755
rect 5946 9679 6054 9755
rect 6426 9679 6534 9755
rect 7194 9679 7302 9755
rect 7674 9679 7782 9755
rect 8442 9679 8550 9755
rect 8922 9679 9030 9755
rect 9690 9679 9798 9755
rect 10170 9679 10278 9755
rect 10938 9679 11046 9755
rect 11418 9679 11526 9755
rect 12186 9679 12294 9755
rect 12666 9679 12774 9755
rect 13434 9679 13542 9755
rect 13914 9679 14022 9755
rect 14682 9679 14790 9755
rect 15162 9679 15270 9755
rect 15930 9679 16038 9755
rect 16410 9679 16518 9755
rect 17178 9679 17286 9755
rect 17658 9679 17766 9755
rect 18426 9679 18534 9755
rect 18906 9679 19014 9755
rect 19674 9679 19782 9755
rect 0 9583 19968 9631
rect 186 9425 294 9535
rect 954 9425 1062 9535
rect 1434 9425 1542 9535
rect 2202 9425 2310 9535
rect 2682 9425 2790 9535
rect 3450 9425 3558 9535
rect 3930 9425 4038 9535
rect 4698 9425 4806 9535
rect 5178 9425 5286 9535
rect 5946 9425 6054 9535
rect 6426 9425 6534 9535
rect 7194 9425 7302 9535
rect 7674 9425 7782 9535
rect 8442 9425 8550 9535
rect 8922 9425 9030 9535
rect 9690 9425 9798 9535
rect 10170 9425 10278 9535
rect 10938 9425 11046 9535
rect 11418 9425 11526 9535
rect 12186 9425 12294 9535
rect 12666 9425 12774 9535
rect 13434 9425 13542 9535
rect 13914 9425 14022 9535
rect 14682 9425 14790 9535
rect 15162 9425 15270 9535
rect 15930 9425 16038 9535
rect 16410 9425 16518 9535
rect 17178 9425 17286 9535
rect 17658 9425 17766 9535
rect 18426 9425 18534 9535
rect 18906 9425 19014 9535
rect 19674 9425 19782 9535
rect 0 9329 19968 9377
rect 186 9205 294 9281
rect 954 9205 1062 9281
rect 1434 9205 1542 9281
rect 2202 9205 2310 9281
rect 2682 9205 2790 9281
rect 3450 9205 3558 9281
rect 3930 9205 4038 9281
rect 4698 9205 4806 9281
rect 5178 9205 5286 9281
rect 5946 9205 6054 9281
rect 6426 9205 6534 9281
rect 7194 9205 7302 9281
rect 7674 9205 7782 9281
rect 8442 9205 8550 9281
rect 8922 9205 9030 9281
rect 9690 9205 9798 9281
rect 10170 9205 10278 9281
rect 10938 9205 11046 9281
rect 11418 9205 11526 9281
rect 12186 9205 12294 9281
rect 12666 9205 12774 9281
rect 13434 9205 13542 9281
rect 13914 9205 14022 9281
rect 14682 9205 14790 9281
rect 15162 9205 15270 9281
rect 15930 9205 16038 9281
rect 16410 9205 16518 9281
rect 17178 9205 17286 9281
rect 17658 9205 17766 9281
rect 18426 9205 18534 9281
rect 18906 9205 19014 9281
rect 19674 9205 19782 9281
rect 0 9109 19968 9157
rect 0 9013 19968 9061
rect 186 8889 294 8965
rect 954 8889 1062 8965
rect 1434 8889 1542 8965
rect 2202 8889 2310 8965
rect 2682 8889 2790 8965
rect 3450 8889 3558 8965
rect 3930 8889 4038 8965
rect 4698 8889 4806 8965
rect 5178 8889 5286 8965
rect 5946 8889 6054 8965
rect 6426 8889 6534 8965
rect 7194 8889 7302 8965
rect 7674 8889 7782 8965
rect 8442 8889 8550 8965
rect 8922 8889 9030 8965
rect 9690 8889 9798 8965
rect 10170 8889 10278 8965
rect 10938 8889 11046 8965
rect 11418 8889 11526 8965
rect 12186 8889 12294 8965
rect 12666 8889 12774 8965
rect 13434 8889 13542 8965
rect 13914 8889 14022 8965
rect 14682 8889 14790 8965
rect 15162 8889 15270 8965
rect 15930 8889 16038 8965
rect 16410 8889 16518 8965
rect 17178 8889 17286 8965
rect 17658 8889 17766 8965
rect 18426 8889 18534 8965
rect 18906 8889 19014 8965
rect 19674 8889 19782 8965
rect 0 8793 19968 8841
rect 186 8635 294 8745
rect 954 8635 1062 8745
rect 1434 8635 1542 8745
rect 2202 8635 2310 8745
rect 2682 8635 2790 8745
rect 3450 8635 3558 8745
rect 3930 8635 4038 8745
rect 4698 8635 4806 8745
rect 5178 8635 5286 8745
rect 5946 8635 6054 8745
rect 6426 8635 6534 8745
rect 7194 8635 7302 8745
rect 7674 8635 7782 8745
rect 8442 8635 8550 8745
rect 8922 8635 9030 8745
rect 9690 8635 9798 8745
rect 10170 8635 10278 8745
rect 10938 8635 11046 8745
rect 11418 8635 11526 8745
rect 12186 8635 12294 8745
rect 12666 8635 12774 8745
rect 13434 8635 13542 8745
rect 13914 8635 14022 8745
rect 14682 8635 14790 8745
rect 15162 8635 15270 8745
rect 15930 8635 16038 8745
rect 16410 8635 16518 8745
rect 17178 8635 17286 8745
rect 17658 8635 17766 8745
rect 18426 8635 18534 8745
rect 18906 8635 19014 8745
rect 19674 8635 19782 8745
rect 0 8539 19968 8587
rect 186 8415 294 8491
rect 954 8415 1062 8491
rect 1434 8415 1542 8491
rect 2202 8415 2310 8491
rect 2682 8415 2790 8491
rect 3450 8415 3558 8491
rect 3930 8415 4038 8491
rect 4698 8415 4806 8491
rect 5178 8415 5286 8491
rect 5946 8415 6054 8491
rect 6426 8415 6534 8491
rect 7194 8415 7302 8491
rect 7674 8415 7782 8491
rect 8442 8415 8550 8491
rect 8922 8415 9030 8491
rect 9690 8415 9798 8491
rect 10170 8415 10278 8491
rect 10938 8415 11046 8491
rect 11418 8415 11526 8491
rect 12186 8415 12294 8491
rect 12666 8415 12774 8491
rect 13434 8415 13542 8491
rect 13914 8415 14022 8491
rect 14682 8415 14790 8491
rect 15162 8415 15270 8491
rect 15930 8415 16038 8491
rect 16410 8415 16518 8491
rect 17178 8415 17286 8491
rect 17658 8415 17766 8491
rect 18426 8415 18534 8491
rect 18906 8415 19014 8491
rect 19674 8415 19782 8491
rect 0 8319 19968 8367
rect 0 8223 19968 8271
rect 186 8099 294 8175
rect 954 8099 1062 8175
rect 1434 8099 1542 8175
rect 2202 8099 2310 8175
rect 2682 8099 2790 8175
rect 3450 8099 3558 8175
rect 3930 8099 4038 8175
rect 4698 8099 4806 8175
rect 5178 8099 5286 8175
rect 5946 8099 6054 8175
rect 6426 8099 6534 8175
rect 7194 8099 7302 8175
rect 7674 8099 7782 8175
rect 8442 8099 8550 8175
rect 8922 8099 9030 8175
rect 9690 8099 9798 8175
rect 10170 8099 10278 8175
rect 10938 8099 11046 8175
rect 11418 8099 11526 8175
rect 12186 8099 12294 8175
rect 12666 8099 12774 8175
rect 13434 8099 13542 8175
rect 13914 8099 14022 8175
rect 14682 8099 14790 8175
rect 15162 8099 15270 8175
rect 15930 8099 16038 8175
rect 16410 8099 16518 8175
rect 17178 8099 17286 8175
rect 17658 8099 17766 8175
rect 18426 8099 18534 8175
rect 18906 8099 19014 8175
rect 19674 8099 19782 8175
rect 0 8003 19968 8051
rect 186 7845 294 7955
rect 954 7845 1062 7955
rect 1434 7845 1542 7955
rect 2202 7845 2310 7955
rect 2682 7845 2790 7955
rect 3450 7845 3558 7955
rect 3930 7845 4038 7955
rect 4698 7845 4806 7955
rect 5178 7845 5286 7955
rect 5946 7845 6054 7955
rect 6426 7845 6534 7955
rect 7194 7845 7302 7955
rect 7674 7845 7782 7955
rect 8442 7845 8550 7955
rect 8922 7845 9030 7955
rect 9690 7845 9798 7955
rect 10170 7845 10278 7955
rect 10938 7845 11046 7955
rect 11418 7845 11526 7955
rect 12186 7845 12294 7955
rect 12666 7845 12774 7955
rect 13434 7845 13542 7955
rect 13914 7845 14022 7955
rect 14682 7845 14790 7955
rect 15162 7845 15270 7955
rect 15930 7845 16038 7955
rect 16410 7845 16518 7955
rect 17178 7845 17286 7955
rect 17658 7845 17766 7955
rect 18426 7845 18534 7955
rect 18906 7845 19014 7955
rect 19674 7845 19782 7955
rect 0 7749 19968 7797
rect 186 7625 294 7701
rect 954 7625 1062 7701
rect 1434 7625 1542 7701
rect 2202 7625 2310 7701
rect 2682 7625 2790 7701
rect 3450 7625 3558 7701
rect 3930 7625 4038 7701
rect 4698 7625 4806 7701
rect 5178 7625 5286 7701
rect 5946 7625 6054 7701
rect 6426 7625 6534 7701
rect 7194 7625 7302 7701
rect 7674 7625 7782 7701
rect 8442 7625 8550 7701
rect 8922 7625 9030 7701
rect 9690 7625 9798 7701
rect 10170 7625 10278 7701
rect 10938 7625 11046 7701
rect 11418 7625 11526 7701
rect 12186 7625 12294 7701
rect 12666 7625 12774 7701
rect 13434 7625 13542 7701
rect 13914 7625 14022 7701
rect 14682 7625 14790 7701
rect 15162 7625 15270 7701
rect 15930 7625 16038 7701
rect 16410 7625 16518 7701
rect 17178 7625 17286 7701
rect 17658 7625 17766 7701
rect 18426 7625 18534 7701
rect 18906 7625 19014 7701
rect 19674 7625 19782 7701
rect 0 7529 19968 7577
rect 0 7433 19968 7481
rect 186 7309 294 7385
rect 954 7309 1062 7385
rect 1434 7309 1542 7385
rect 2202 7309 2310 7385
rect 2682 7309 2790 7385
rect 3450 7309 3558 7385
rect 3930 7309 4038 7385
rect 4698 7309 4806 7385
rect 5178 7309 5286 7385
rect 5946 7309 6054 7385
rect 6426 7309 6534 7385
rect 7194 7309 7302 7385
rect 7674 7309 7782 7385
rect 8442 7309 8550 7385
rect 8922 7309 9030 7385
rect 9690 7309 9798 7385
rect 10170 7309 10278 7385
rect 10938 7309 11046 7385
rect 11418 7309 11526 7385
rect 12186 7309 12294 7385
rect 12666 7309 12774 7385
rect 13434 7309 13542 7385
rect 13914 7309 14022 7385
rect 14682 7309 14790 7385
rect 15162 7309 15270 7385
rect 15930 7309 16038 7385
rect 16410 7309 16518 7385
rect 17178 7309 17286 7385
rect 17658 7309 17766 7385
rect 18426 7309 18534 7385
rect 18906 7309 19014 7385
rect 19674 7309 19782 7385
rect 0 7213 19968 7261
rect 186 7055 294 7165
rect 954 7055 1062 7165
rect 1434 7055 1542 7165
rect 2202 7055 2310 7165
rect 2682 7055 2790 7165
rect 3450 7055 3558 7165
rect 3930 7055 4038 7165
rect 4698 7055 4806 7165
rect 5178 7055 5286 7165
rect 5946 7055 6054 7165
rect 6426 7055 6534 7165
rect 7194 7055 7302 7165
rect 7674 7055 7782 7165
rect 8442 7055 8550 7165
rect 8922 7055 9030 7165
rect 9690 7055 9798 7165
rect 10170 7055 10278 7165
rect 10938 7055 11046 7165
rect 11418 7055 11526 7165
rect 12186 7055 12294 7165
rect 12666 7055 12774 7165
rect 13434 7055 13542 7165
rect 13914 7055 14022 7165
rect 14682 7055 14790 7165
rect 15162 7055 15270 7165
rect 15930 7055 16038 7165
rect 16410 7055 16518 7165
rect 17178 7055 17286 7165
rect 17658 7055 17766 7165
rect 18426 7055 18534 7165
rect 18906 7055 19014 7165
rect 19674 7055 19782 7165
rect 0 6959 19968 7007
rect 186 6835 294 6911
rect 954 6835 1062 6911
rect 1434 6835 1542 6911
rect 2202 6835 2310 6911
rect 2682 6835 2790 6911
rect 3450 6835 3558 6911
rect 3930 6835 4038 6911
rect 4698 6835 4806 6911
rect 5178 6835 5286 6911
rect 5946 6835 6054 6911
rect 6426 6835 6534 6911
rect 7194 6835 7302 6911
rect 7674 6835 7782 6911
rect 8442 6835 8550 6911
rect 8922 6835 9030 6911
rect 9690 6835 9798 6911
rect 10170 6835 10278 6911
rect 10938 6835 11046 6911
rect 11418 6835 11526 6911
rect 12186 6835 12294 6911
rect 12666 6835 12774 6911
rect 13434 6835 13542 6911
rect 13914 6835 14022 6911
rect 14682 6835 14790 6911
rect 15162 6835 15270 6911
rect 15930 6835 16038 6911
rect 16410 6835 16518 6911
rect 17178 6835 17286 6911
rect 17658 6835 17766 6911
rect 18426 6835 18534 6911
rect 18906 6835 19014 6911
rect 19674 6835 19782 6911
rect 0 6739 19968 6787
rect 0 6643 19968 6691
rect 186 6519 294 6595
rect 954 6519 1062 6595
rect 1434 6519 1542 6595
rect 2202 6519 2310 6595
rect 2682 6519 2790 6595
rect 3450 6519 3558 6595
rect 3930 6519 4038 6595
rect 4698 6519 4806 6595
rect 5178 6519 5286 6595
rect 5946 6519 6054 6595
rect 6426 6519 6534 6595
rect 7194 6519 7302 6595
rect 7674 6519 7782 6595
rect 8442 6519 8550 6595
rect 8922 6519 9030 6595
rect 9690 6519 9798 6595
rect 10170 6519 10278 6595
rect 10938 6519 11046 6595
rect 11418 6519 11526 6595
rect 12186 6519 12294 6595
rect 12666 6519 12774 6595
rect 13434 6519 13542 6595
rect 13914 6519 14022 6595
rect 14682 6519 14790 6595
rect 15162 6519 15270 6595
rect 15930 6519 16038 6595
rect 16410 6519 16518 6595
rect 17178 6519 17286 6595
rect 17658 6519 17766 6595
rect 18426 6519 18534 6595
rect 18906 6519 19014 6595
rect 19674 6519 19782 6595
rect 0 6423 19968 6471
rect 186 6265 294 6375
rect 954 6265 1062 6375
rect 1434 6265 1542 6375
rect 2202 6265 2310 6375
rect 2682 6265 2790 6375
rect 3450 6265 3558 6375
rect 3930 6265 4038 6375
rect 4698 6265 4806 6375
rect 5178 6265 5286 6375
rect 5946 6265 6054 6375
rect 6426 6265 6534 6375
rect 7194 6265 7302 6375
rect 7674 6265 7782 6375
rect 8442 6265 8550 6375
rect 8922 6265 9030 6375
rect 9690 6265 9798 6375
rect 10170 6265 10278 6375
rect 10938 6265 11046 6375
rect 11418 6265 11526 6375
rect 12186 6265 12294 6375
rect 12666 6265 12774 6375
rect 13434 6265 13542 6375
rect 13914 6265 14022 6375
rect 14682 6265 14790 6375
rect 15162 6265 15270 6375
rect 15930 6265 16038 6375
rect 16410 6265 16518 6375
rect 17178 6265 17286 6375
rect 17658 6265 17766 6375
rect 18426 6265 18534 6375
rect 18906 6265 19014 6375
rect 19674 6265 19782 6375
rect 0 6169 19968 6217
rect 186 6045 294 6121
rect 954 6045 1062 6121
rect 1434 6045 1542 6121
rect 2202 6045 2310 6121
rect 2682 6045 2790 6121
rect 3450 6045 3558 6121
rect 3930 6045 4038 6121
rect 4698 6045 4806 6121
rect 5178 6045 5286 6121
rect 5946 6045 6054 6121
rect 6426 6045 6534 6121
rect 7194 6045 7302 6121
rect 7674 6045 7782 6121
rect 8442 6045 8550 6121
rect 8922 6045 9030 6121
rect 9690 6045 9798 6121
rect 10170 6045 10278 6121
rect 10938 6045 11046 6121
rect 11418 6045 11526 6121
rect 12186 6045 12294 6121
rect 12666 6045 12774 6121
rect 13434 6045 13542 6121
rect 13914 6045 14022 6121
rect 14682 6045 14790 6121
rect 15162 6045 15270 6121
rect 15930 6045 16038 6121
rect 16410 6045 16518 6121
rect 17178 6045 17286 6121
rect 17658 6045 17766 6121
rect 18426 6045 18534 6121
rect 18906 6045 19014 6121
rect 19674 6045 19782 6121
rect 0 5949 19968 5997
rect 0 5853 19968 5901
rect 186 5729 294 5805
rect 954 5729 1062 5805
rect 1434 5729 1542 5805
rect 2202 5729 2310 5805
rect 2682 5729 2790 5805
rect 3450 5729 3558 5805
rect 3930 5729 4038 5805
rect 4698 5729 4806 5805
rect 5178 5729 5286 5805
rect 5946 5729 6054 5805
rect 6426 5729 6534 5805
rect 7194 5729 7302 5805
rect 7674 5729 7782 5805
rect 8442 5729 8550 5805
rect 8922 5729 9030 5805
rect 9690 5729 9798 5805
rect 10170 5729 10278 5805
rect 10938 5729 11046 5805
rect 11418 5729 11526 5805
rect 12186 5729 12294 5805
rect 12666 5729 12774 5805
rect 13434 5729 13542 5805
rect 13914 5729 14022 5805
rect 14682 5729 14790 5805
rect 15162 5729 15270 5805
rect 15930 5729 16038 5805
rect 16410 5729 16518 5805
rect 17178 5729 17286 5805
rect 17658 5729 17766 5805
rect 18426 5729 18534 5805
rect 18906 5729 19014 5805
rect 19674 5729 19782 5805
rect 0 5633 19968 5681
rect 186 5475 294 5585
rect 954 5475 1062 5585
rect 1434 5475 1542 5585
rect 2202 5475 2310 5585
rect 2682 5475 2790 5585
rect 3450 5475 3558 5585
rect 3930 5475 4038 5585
rect 4698 5475 4806 5585
rect 5178 5475 5286 5585
rect 5946 5475 6054 5585
rect 6426 5475 6534 5585
rect 7194 5475 7302 5585
rect 7674 5475 7782 5585
rect 8442 5475 8550 5585
rect 8922 5475 9030 5585
rect 9690 5475 9798 5585
rect 10170 5475 10278 5585
rect 10938 5475 11046 5585
rect 11418 5475 11526 5585
rect 12186 5475 12294 5585
rect 12666 5475 12774 5585
rect 13434 5475 13542 5585
rect 13914 5475 14022 5585
rect 14682 5475 14790 5585
rect 15162 5475 15270 5585
rect 15930 5475 16038 5585
rect 16410 5475 16518 5585
rect 17178 5475 17286 5585
rect 17658 5475 17766 5585
rect 18426 5475 18534 5585
rect 18906 5475 19014 5585
rect 19674 5475 19782 5585
rect 0 5379 19968 5427
rect 186 5255 294 5331
rect 954 5255 1062 5331
rect 1434 5255 1542 5331
rect 2202 5255 2310 5331
rect 2682 5255 2790 5331
rect 3450 5255 3558 5331
rect 3930 5255 4038 5331
rect 4698 5255 4806 5331
rect 5178 5255 5286 5331
rect 5946 5255 6054 5331
rect 6426 5255 6534 5331
rect 7194 5255 7302 5331
rect 7674 5255 7782 5331
rect 8442 5255 8550 5331
rect 8922 5255 9030 5331
rect 9690 5255 9798 5331
rect 10170 5255 10278 5331
rect 10938 5255 11046 5331
rect 11418 5255 11526 5331
rect 12186 5255 12294 5331
rect 12666 5255 12774 5331
rect 13434 5255 13542 5331
rect 13914 5255 14022 5331
rect 14682 5255 14790 5331
rect 15162 5255 15270 5331
rect 15930 5255 16038 5331
rect 16410 5255 16518 5331
rect 17178 5255 17286 5331
rect 17658 5255 17766 5331
rect 18426 5255 18534 5331
rect 18906 5255 19014 5331
rect 19674 5255 19782 5331
rect 0 5159 19968 5207
rect 0 5063 19968 5111
rect 186 4939 294 5015
rect 954 4939 1062 5015
rect 1434 4939 1542 5015
rect 2202 4939 2310 5015
rect 2682 4939 2790 5015
rect 3450 4939 3558 5015
rect 3930 4939 4038 5015
rect 4698 4939 4806 5015
rect 5178 4939 5286 5015
rect 5946 4939 6054 5015
rect 6426 4939 6534 5015
rect 7194 4939 7302 5015
rect 7674 4939 7782 5015
rect 8442 4939 8550 5015
rect 8922 4939 9030 5015
rect 9690 4939 9798 5015
rect 10170 4939 10278 5015
rect 10938 4939 11046 5015
rect 11418 4939 11526 5015
rect 12186 4939 12294 5015
rect 12666 4939 12774 5015
rect 13434 4939 13542 5015
rect 13914 4939 14022 5015
rect 14682 4939 14790 5015
rect 15162 4939 15270 5015
rect 15930 4939 16038 5015
rect 16410 4939 16518 5015
rect 17178 4939 17286 5015
rect 17658 4939 17766 5015
rect 18426 4939 18534 5015
rect 18906 4939 19014 5015
rect 19674 4939 19782 5015
rect 0 4843 19968 4891
rect 186 4685 294 4795
rect 954 4685 1062 4795
rect 1434 4685 1542 4795
rect 2202 4685 2310 4795
rect 2682 4685 2790 4795
rect 3450 4685 3558 4795
rect 3930 4685 4038 4795
rect 4698 4685 4806 4795
rect 5178 4685 5286 4795
rect 5946 4685 6054 4795
rect 6426 4685 6534 4795
rect 7194 4685 7302 4795
rect 7674 4685 7782 4795
rect 8442 4685 8550 4795
rect 8922 4685 9030 4795
rect 9690 4685 9798 4795
rect 10170 4685 10278 4795
rect 10938 4685 11046 4795
rect 11418 4685 11526 4795
rect 12186 4685 12294 4795
rect 12666 4685 12774 4795
rect 13434 4685 13542 4795
rect 13914 4685 14022 4795
rect 14682 4685 14790 4795
rect 15162 4685 15270 4795
rect 15930 4685 16038 4795
rect 16410 4685 16518 4795
rect 17178 4685 17286 4795
rect 17658 4685 17766 4795
rect 18426 4685 18534 4795
rect 18906 4685 19014 4795
rect 19674 4685 19782 4795
rect 0 4589 19968 4637
rect 186 4465 294 4541
rect 954 4465 1062 4541
rect 1434 4465 1542 4541
rect 2202 4465 2310 4541
rect 2682 4465 2790 4541
rect 3450 4465 3558 4541
rect 3930 4465 4038 4541
rect 4698 4465 4806 4541
rect 5178 4465 5286 4541
rect 5946 4465 6054 4541
rect 6426 4465 6534 4541
rect 7194 4465 7302 4541
rect 7674 4465 7782 4541
rect 8442 4465 8550 4541
rect 8922 4465 9030 4541
rect 9690 4465 9798 4541
rect 10170 4465 10278 4541
rect 10938 4465 11046 4541
rect 11418 4465 11526 4541
rect 12186 4465 12294 4541
rect 12666 4465 12774 4541
rect 13434 4465 13542 4541
rect 13914 4465 14022 4541
rect 14682 4465 14790 4541
rect 15162 4465 15270 4541
rect 15930 4465 16038 4541
rect 16410 4465 16518 4541
rect 17178 4465 17286 4541
rect 17658 4465 17766 4541
rect 18426 4465 18534 4541
rect 18906 4465 19014 4541
rect 19674 4465 19782 4541
rect 0 4369 19968 4417
rect 0 4273 19968 4321
rect 186 4149 294 4225
rect 954 4149 1062 4225
rect 1434 4149 1542 4225
rect 2202 4149 2310 4225
rect 2682 4149 2790 4225
rect 3450 4149 3558 4225
rect 3930 4149 4038 4225
rect 4698 4149 4806 4225
rect 5178 4149 5286 4225
rect 5946 4149 6054 4225
rect 6426 4149 6534 4225
rect 7194 4149 7302 4225
rect 7674 4149 7782 4225
rect 8442 4149 8550 4225
rect 8922 4149 9030 4225
rect 9690 4149 9798 4225
rect 10170 4149 10278 4225
rect 10938 4149 11046 4225
rect 11418 4149 11526 4225
rect 12186 4149 12294 4225
rect 12666 4149 12774 4225
rect 13434 4149 13542 4225
rect 13914 4149 14022 4225
rect 14682 4149 14790 4225
rect 15162 4149 15270 4225
rect 15930 4149 16038 4225
rect 16410 4149 16518 4225
rect 17178 4149 17286 4225
rect 17658 4149 17766 4225
rect 18426 4149 18534 4225
rect 18906 4149 19014 4225
rect 19674 4149 19782 4225
rect 0 4053 19968 4101
rect 186 3895 294 4005
rect 954 3895 1062 4005
rect 1434 3895 1542 4005
rect 2202 3895 2310 4005
rect 2682 3895 2790 4005
rect 3450 3895 3558 4005
rect 3930 3895 4038 4005
rect 4698 3895 4806 4005
rect 5178 3895 5286 4005
rect 5946 3895 6054 4005
rect 6426 3895 6534 4005
rect 7194 3895 7302 4005
rect 7674 3895 7782 4005
rect 8442 3895 8550 4005
rect 8922 3895 9030 4005
rect 9690 3895 9798 4005
rect 10170 3895 10278 4005
rect 10938 3895 11046 4005
rect 11418 3895 11526 4005
rect 12186 3895 12294 4005
rect 12666 3895 12774 4005
rect 13434 3895 13542 4005
rect 13914 3895 14022 4005
rect 14682 3895 14790 4005
rect 15162 3895 15270 4005
rect 15930 3895 16038 4005
rect 16410 3895 16518 4005
rect 17178 3895 17286 4005
rect 17658 3895 17766 4005
rect 18426 3895 18534 4005
rect 18906 3895 19014 4005
rect 19674 3895 19782 4005
rect 0 3799 19968 3847
rect 186 3675 294 3751
rect 954 3675 1062 3751
rect 1434 3675 1542 3751
rect 2202 3675 2310 3751
rect 2682 3675 2790 3751
rect 3450 3675 3558 3751
rect 3930 3675 4038 3751
rect 4698 3675 4806 3751
rect 5178 3675 5286 3751
rect 5946 3675 6054 3751
rect 6426 3675 6534 3751
rect 7194 3675 7302 3751
rect 7674 3675 7782 3751
rect 8442 3675 8550 3751
rect 8922 3675 9030 3751
rect 9690 3675 9798 3751
rect 10170 3675 10278 3751
rect 10938 3675 11046 3751
rect 11418 3675 11526 3751
rect 12186 3675 12294 3751
rect 12666 3675 12774 3751
rect 13434 3675 13542 3751
rect 13914 3675 14022 3751
rect 14682 3675 14790 3751
rect 15162 3675 15270 3751
rect 15930 3675 16038 3751
rect 16410 3675 16518 3751
rect 17178 3675 17286 3751
rect 17658 3675 17766 3751
rect 18426 3675 18534 3751
rect 18906 3675 19014 3751
rect 19674 3675 19782 3751
rect 0 3579 19968 3627
rect 0 3483 19968 3531
rect 186 3359 294 3435
rect 954 3359 1062 3435
rect 1434 3359 1542 3435
rect 2202 3359 2310 3435
rect 2682 3359 2790 3435
rect 3450 3359 3558 3435
rect 3930 3359 4038 3435
rect 4698 3359 4806 3435
rect 5178 3359 5286 3435
rect 5946 3359 6054 3435
rect 6426 3359 6534 3435
rect 7194 3359 7302 3435
rect 7674 3359 7782 3435
rect 8442 3359 8550 3435
rect 8922 3359 9030 3435
rect 9690 3359 9798 3435
rect 10170 3359 10278 3435
rect 10938 3359 11046 3435
rect 11418 3359 11526 3435
rect 12186 3359 12294 3435
rect 12666 3359 12774 3435
rect 13434 3359 13542 3435
rect 13914 3359 14022 3435
rect 14682 3359 14790 3435
rect 15162 3359 15270 3435
rect 15930 3359 16038 3435
rect 16410 3359 16518 3435
rect 17178 3359 17286 3435
rect 17658 3359 17766 3435
rect 18426 3359 18534 3435
rect 18906 3359 19014 3435
rect 19674 3359 19782 3435
rect 0 3263 19968 3311
rect 186 3105 294 3215
rect 954 3105 1062 3215
rect 1434 3105 1542 3215
rect 2202 3105 2310 3215
rect 2682 3105 2790 3215
rect 3450 3105 3558 3215
rect 3930 3105 4038 3215
rect 4698 3105 4806 3215
rect 5178 3105 5286 3215
rect 5946 3105 6054 3215
rect 6426 3105 6534 3215
rect 7194 3105 7302 3215
rect 7674 3105 7782 3215
rect 8442 3105 8550 3215
rect 8922 3105 9030 3215
rect 9690 3105 9798 3215
rect 10170 3105 10278 3215
rect 10938 3105 11046 3215
rect 11418 3105 11526 3215
rect 12186 3105 12294 3215
rect 12666 3105 12774 3215
rect 13434 3105 13542 3215
rect 13914 3105 14022 3215
rect 14682 3105 14790 3215
rect 15162 3105 15270 3215
rect 15930 3105 16038 3215
rect 16410 3105 16518 3215
rect 17178 3105 17286 3215
rect 17658 3105 17766 3215
rect 18426 3105 18534 3215
rect 18906 3105 19014 3215
rect 19674 3105 19782 3215
rect 0 3009 19968 3057
rect 186 2885 294 2961
rect 954 2885 1062 2961
rect 1434 2885 1542 2961
rect 2202 2885 2310 2961
rect 2682 2885 2790 2961
rect 3450 2885 3558 2961
rect 3930 2885 4038 2961
rect 4698 2885 4806 2961
rect 5178 2885 5286 2961
rect 5946 2885 6054 2961
rect 6426 2885 6534 2961
rect 7194 2885 7302 2961
rect 7674 2885 7782 2961
rect 8442 2885 8550 2961
rect 8922 2885 9030 2961
rect 9690 2885 9798 2961
rect 10170 2885 10278 2961
rect 10938 2885 11046 2961
rect 11418 2885 11526 2961
rect 12186 2885 12294 2961
rect 12666 2885 12774 2961
rect 13434 2885 13542 2961
rect 13914 2885 14022 2961
rect 14682 2885 14790 2961
rect 15162 2885 15270 2961
rect 15930 2885 16038 2961
rect 16410 2885 16518 2961
rect 17178 2885 17286 2961
rect 17658 2885 17766 2961
rect 18426 2885 18534 2961
rect 18906 2885 19014 2961
rect 19674 2885 19782 2961
rect 0 2789 19968 2837
rect 0 2693 19968 2741
rect 186 2569 294 2645
rect 954 2569 1062 2645
rect 1434 2569 1542 2645
rect 2202 2569 2310 2645
rect 2682 2569 2790 2645
rect 3450 2569 3558 2645
rect 3930 2569 4038 2645
rect 4698 2569 4806 2645
rect 5178 2569 5286 2645
rect 5946 2569 6054 2645
rect 6426 2569 6534 2645
rect 7194 2569 7302 2645
rect 7674 2569 7782 2645
rect 8442 2569 8550 2645
rect 8922 2569 9030 2645
rect 9690 2569 9798 2645
rect 10170 2569 10278 2645
rect 10938 2569 11046 2645
rect 11418 2569 11526 2645
rect 12186 2569 12294 2645
rect 12666 2569 12774 2645
rect 13434 2569 13542 2645
rect 13914 2569 14022 2645
rect 14682 2569 14790 2645
rect 15162 2569 15270 2645
rect 15930 2569 16038 2645
rect 16410 2569 16518 2645
rect 17178 2569 17286 2645
rect 17658 2569 17766 2645
rect 18426 2569 18534 2645
rect 18906 2569 19014 2645
rect 19674 2569 19782 2645
rect 0 2473 19968 2521
rect 186 2315 294 2425
rect 954 2315 1062 2425
rect 1434 2315 1542 2425
rect 2202 2315 2310 2425
rect 2682 2315 2790 2425
rect 3450 2315 3558 2425
rect 3930 2315 4038 2425
rect 4698 2315 4806 2425
rect 5178 2315 5286 2425
rect 5946 2315 6054 2425
rect 6426 2315 6534 2425
rect 7194 2315 7302 2425
rect 7674 2315 7782 2425
rect 8442 2315 8550 2425
rect 8922 2315 9030 2425
rect 9690 2315 9798 2425
rect 10170 2315 10278 2425
rect 10938 2315 11046 2425
rect 11418 2315 11526 2425
rect 12186 2315 12294 2425
rect 12666 2315 12774 2425
rect 13434 2315 13542 2425
rect 13914 2315 14022 2425
rect 14682 2315 14790 2425
rect 15162 2315 15270 2425
rect 15930 2315 16038 2425
rect 16410 2315 16518 2425
rect 17178 2315 17286 2425
rect 17658 2315 17766 2425
rect 18426 2315 18534 2425
rect 18906 2315 19014 2425
rect 19674 2315 19782 2425
rect 0 2219 19968 2267
rect 186 2095 294 2171
rect 954 2095 1062 2171
rect 1434 2095 1542 2171
rect 2202 2095 2310 2171
rect 2682 2095 2790 2171
rect 3450 2095 3558 2171
rect 3930 2095 4038 2171
rect 4698 2095 4806 2171
rect 5178 2095 5286 2171
rect 5946 2095 6054 2171
rect 6426 2095 6534 2171
rect 7194 2095 7302 2171
rect 7674 2095 7782 2171
rect 8442 2095 8550 2171
rect 8922 2095 9030 2171
rect 9690 2095 9798 2171
rect 10170 2095 10278 2171
rect 10938 2095 11046 2171
rect 11418 2095 11526 2171
rect 12186 2095 12294 2171
rect 12666 2095 12774 2171
rect 13434 2095 13542 2171
rect 13914 2095 14022 2171
rect 14682 2095 14790 2171
rect 15162 2095 15270 2171
rect 15930 2095 16038 2171
rect 16410 2095 16518 2171
rect 17178 2095 17286 2171
rect 17658 2095 17766 2171
rect 18426 2095 18534 2171
rect 18906 2095 19014 2171
rect 19674 2095 19782 2171
rect 0 1999 19968 2047
rect 0 1903 19968 1951
rect 186 1779 294 1855
rect 954 1779 1062 1855
rect 1434 1779 1542 1855
rect 2202 1779 2310 1855
rect 2682 1779 2790 1855
rect 3450 1779 3558 1855
rect 3930 1779 4038 1855
rect 4698 1779 4806 1855
rect 5178 1779 5286 1855
rect 5946 1779 6054 1855
rect 6426 1779 6534 1855
rect 7194 1779 7302 1855
rect 7674 1779 7782 1855
rect 8442 1779 8550 1855
rect 8922 1779 9030 1855
rect 9690 1779 9798 1855
rect 10170 1779 10278 1855
rect 10938 1779 11046 1855
rect 11418 1779 11526 1855
rect 12186 1779 12294 1855
rect 12666 1779 12774 1855
rect 13434 1779 13542 1855
rect 13914 1779 14022 1855
rect 14682 1779 14790 1855
rect 15162 1779 15270 1855
rect 15930 1779 16038 1855
rect 16410 1779 16518 1855
rect 17178 1779 17286 1855
rect 17658 1779 17766 1855
rect 18426 1779 18534 1855
rect 18906 1779 19014 1855
rect 19674 1779 19782 1855
rect 0 1683 19968 1731
rect 186 1525 294 1635
rect 954 1525 1062 1635
rect 1434 1525 1542 1635
rect 2202 1525 2310 1635
rect 2682 1525 2790 1635
rect 3450 1525 3558 1635
rect 3930 1525 4038 1635
rect 4698 1525 4806 1635
rect 5178 1525 5286 1635
rect 5946 1525 6054 1635
rect 6426 1525 6534 1635
rect 7194 1525 7302 1635
rect 7674 1525 7782 1635
rect 8442 1525 8550 1635
rect 8922 1525 9030 1635
rect 9690 1525 9798 1635
rect 10170 1525 10278 1635
rect 10938 1525 11046 1635
rect 11418 1525 11526 1635
rect 12186 1525 12294 1635
rect 12666 1525 12774 1635
rect 13434 1525 13542 1635
rect 13914 1525 14022 1635
rect 14682 1525 14790 1635
rect 15162 1525 15270 1635
rect 15930 1525 16038 1635
rect 16410 1525 16518 1635
rect 17178 1525 17286 1635
rect 17658 1525 17766 1635
rect 18426 1525 18534 1635
rect 18906 1525 19014 1635
rect 19674 1525 19782 1635
rect 0 1429 19968 1477
rect 186 1305 294 1381
rect 954 1305 1062 1381
rect 1434 1305 1542 1381
rect 2202 1305 2310 1381
rect 2682 1305 2790 1381
rect 3450 1305 3558 1381
rect 3930 1305 4038 1381
rect 4698 1305 4806 1381
rect 5178 1305 5286 1381
rect 5946 1305 6054 1381
rect 6426 1305 6534 1381
rect 7194 1305 7302 1381
rect 7674 1305 7782 1381
rect 8442 1305 8550 1381
rect 8922 1305 9030 1381
rect 9690 1305 9798 1381
rect 10170 1305 10278 1381
rect 10938 1305 11046 1381
rect 11418 1305 11526 1381
rect 12186 1305 12294 1381
rect 12666 1305 12774 1381
rect 13434 1305 13542 1381
rect 13914 1305 14022 1381
rect 14682 1305 14790 1381
rect 15162 1305 15270 1381
rect 15930 1305 16038 1381
rect 16410 1305 16518 1381
rect 17178 1305 17286 1381
rect 17658 1305 17766 1381
rect 18426 1305 18534 1381
rect 18906 1305 19014 1381
rect 19674 1305 19782 1381
rect 0 1209 19968 1257
rect 0 1113 19968 1161
rect 186 989 294 1065
rect 954 989 1062 1065
rect 1434 989 1542 1065
rect 2202 989 2310 1065
rect 2682 989 2790 1065
rect 3450 989 3558 1065
rect 3930 989 4038 1065
rect 4698 989 4806 1065
rect 5178 989 5286 1065
rect 5946 989 6054 1065
rect 6426 989 6534 1065
rect 7194 989 7302 1065
rect 7674 989 7782 1065
rect 8442 989 8550 1065
rect 8922 989 9030 1065
rect 9690 989 9798 1065
rect 10170 989 10278 1065
rect 10938 989 11046 1065
rect 11418 989 11526 1065
rect 12186 989 12294 1065
rect 12666 989 12774 1065
rect 13434 989 13542 1065
rect 13914 989 14022 1065
rect 14682 989 14790 1065
rect 15162 989 15270 1065
rect 15930 989 16038 1065
rect 16410 989 16518 1065
rect 17178 989 17286 1065
rect 17658 989 17766 1065
rect 18426 989 18534 1065
rect 18906 989 19014 1065
rect 19674 989 19782 1065
rect 0 893 19968 941
rect 186 735 294 845
rect 954 735 1062 845
rect 1434 735 1542 845
rect 2202 735 2310 845
rect 2682 735 2790 845
rect 3450 735 3558 845
rect 3930 735 4038 845
rect 4698 735 4806 845
rect 5178 735 5286 845
rect 5946 735 6054 845
rect 6426 735 6534 845
rect 7194 735 7302 845
rect 7674 735 7782 845
rect 8442 735 8550 845
rect 8922 735 9030 845
rect 9690 735 9798 845
rect 10170 735 10278 845
rect 10938 735 11046 845
rect 11418 735 11526 845
rect 12186 735 12294 845
rect 12666 735 12774 845
rect 13434 735 13542 845
rect 13914 735 14022 845
rect 14682 735 14790 845
rect 15162 735 15270 845
rect 15930 735 16038 845
rect 16410 735 16518 845
rect 17178 735 17286 845
rect 17658 735 17766 845
rect 18426 735 18534 845
rect 18906 735 19014 845
rect 19674 735 19782 845
rect 0 639 19968 687
rect 186 515 294 591
rect 954 515 1062 591
rect 1434 515 1542 591
rect 2202 515 2310 591
rect 2682 515 2790 591
rect 3450 515 3558 591
rect 3930 515 4038 591
rect 4698 515 4806 591
rect 5178 515 5286 591
rect 5946 515 6054 591
rect 6426 515 6534 591
rect 7194 515 7302 591
rect 7674 515 7782 591
rect 8442 515 8550 591
rect 8922 515 9030 591
rect 9690 515 9798 591
rect 10170 515 10278 591
rect 10938 515 11046 591
rect 11418 515 11526 591
rect 12186 515 12294 591
rect 12666 515 12774 591
rect 13434 515 13542 591
rect 13914 515 14022 591
rect 14682 515 14790 591
rect 15162 515 15270 591
rect 15930 515 16038 591
rect 16410 515 16518 591
rect 17178 515 17286 591
rect 17658 515 17766 591
rect 18426 515 18534 591
rect 18906 515 19014 591
rect 19674 515 19782 591
rect 0 419 19968 467
rect 0 323 19968 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 0 103 19968 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_0
timestamp 1435914306
transform -1 0 19968 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1
timestamp 1435914306
transform -1 0 19968 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2
timestamp 1435914306
transform -1 0 19968 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_3
timestamp 1435914306
transform -1 0 19968 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_4
timestamp 1435914306
transform -1 0 19968 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_5
timestamp 1435914306
transform -1 0 19968 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_6
timestamp 1435914306
transform -1 0 19968 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_7
timestamp 1435914306
transform -1 0 19968 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_8
timestamp 1435914306
transform -1 0 19968 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_9
timestamp 1435914306
transform -1 0 19968 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_10
timestamp 1435914306
transform -1 0 19968 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_11
timestamp 1435914306
transform -1 0 19968 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_12
timestamp 1435914306
transform -1 0 19968 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_13
timestamp 1435914306
transform -1 0 19968 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_14
timestamp 1435914306
transform -1 0 19968 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_15
timestamp 1435914306
transform -1 0 19968 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_16
timestamp 1435914306
transform -1 0 19968 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_17
timestamp 1435914306
transform -1 0 19968 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_18
timestamp 1435914306
transform -1 0 19968 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_19
timestamp 1435914306
transform -1 0 19968 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_20
timestamp 1435914306
transform -1 0 19968 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_21
timestamp 1435914306
transform -1 0 19968 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_22
timestamp 1435914306
transform -1 0 19968 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_23
timestamp 1435914306
transform -1 0 19968 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_24
timestamp 1435914306
transform -1 0 19968 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_25
timestamp 1435914306
transform -1 0 19968 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_26
timestamp 1435914306
transform -1 0 19968 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_27
timestamp 1435914306
transform -1 0 19968 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_28
timestamp 1435914306
transform -1 0 19968 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_29
timestamp 1435914306
transform -1 0 19968 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_30
timestamp 1435914306
transform -1 0 19968 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_31
timestamp 1435914306
transform -1 0 19968 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_32
timestamp 1435914306
transform -1 0 19968 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_33
timestamp 1435914306
transform -1 0 19968 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_34
timestamp 1435914306
transform -1 0 19968 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_35
timestamp 1435914306
transform -1 0 19968 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_36
timestamp 1435914306
transform -1 0 19968 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_37
timestamp 1435914306
transform -1 0 19968 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_38
timestamp 1435914306
transform -1 0 19968 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_39
timestamp 1435914306
transform -1 0 19968 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_40
timestamp 1435914306
transform -1 0 19968 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_41
timestamp 1435914306
transform -1 0 19968 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_42
timestamp 1435914306
transform -1 0 19968 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_43
timestamp 1435914306
transform -1 0 19968 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_44
timestamp 1435914306
transform -1 0 19968 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_45
timestamp 1435914306
transform -1 0 19968 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_46
timestamp 1435914306
transform -1 0 19968 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_47
timestamp 1435914306
transform -1 0 19968 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_48
timestamp 1435914306
transform -1 0 19968 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_49
timestamp 1435914306
transform -1 0 19968 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_50
timestamp 1435914306
transform -1 0 19968 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_51
timestamp 1435914306
transform -1 0 19968 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_52
timestamp 1435914306
transform -1 0 19968 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_53
timestamp 1435914306
transform -1 0 19968 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_54
timestamp 1435914306
transform -1 0 19968 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_55
timestamp 1435914306
transform -1 0 19968 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_56
timestamp 1435914306
transform -1 0 19968 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_57
timestamp 1435914306
transform -1 0 19968 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_58
timestamp 1435914306
transform -1 0 19968 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_59
timestamp 1435914306
transform -1 0 19968 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_60
timestamp 1435914306
transform -1 0 19968 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_61
timestamp 1435914306
transform -1 0 19968 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_62
timestamp 1435914306
transform -1 0 19968 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_63
timestamp 1435914306
transform -1 0 19968 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_64
timestamp 1435914306
transform 1 0 18720 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_65
timestamp 1435914306
transform 1 0 18720 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_66
timestamp 1435914306
transform 1 0 18720 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_67
timestamp 1435914306
transform 1 0 18720 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_68
timestamp 1435914306
transform 1 0 18720 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_69
timestamp 1435914306
transform 1 0 18720 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_70
timestamp 1435914306
transform 1 0 18720 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_71
timestamp 1435914306
transform 1 0 18720 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_72
timestamp 1435914306
transform 1 0 18720 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_73
timestamp 1435914306
transform 1 0 18720 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_74
timestamp 1435914306
transform 1 0 18720 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_75
timestamp 1435914306
transform 1 0 18720 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_76
timestamp 1435914306
transform 1 0 18720 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_77
timestamp 1435914306
transform 1 0 18720 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_78
timestamp 1435914306
transform 1 0 18720 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_79
timestamp 1435914306
transform 1 0 18720 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_80
timestamp 1435914306
transform 1 0 18720 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_81
timestamp 1435914306
transform 1 0 18720 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_82
timestamp 1435914306
transform 1 0 18720 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_83
timestamp 1435914306
transform 1 0 18720 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_84
timestamp 1435914306
transform 1 0 18720 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_85
timestamp 1435914306
transform 1 0 18720 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_86
timestamp 1435914306
transform 1 0 18720 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_87
timestamp 1435914306
transform 1 0 18720 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_88
timestamp 1435914306
transform 1 0 18720 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_89
timestamp 1435914306
transform 1 0 18720 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_90
timestamp 1435914306
transform 1 0 18720 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_91
timestamp 1435914306
transform 1 0 18720 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_92
timestamp 1435914306
transform 1 0 18720 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_93
timestamp 1435914306
transform 1 0 18720 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_94
timestamp 1435914306
transform 1 0 18720 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_95
timestamp 1435914306
transform 1 0 18720 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_96
timestamp 1435914306
transform 1 0 18720 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_97
timestamp 1435914306
transform 1 0 18720 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_98
timestamp 1435914306
transform 1 0 18720 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_99
timestamp 1435914306
transform 1 0 18720 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_100
timestamp 1435914306
transform 1 0 18720 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_101
timestamp 1435914306
transform 1 0 18720 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_102
timestamp 1435914306
transform 1 0 18720 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_103
timestamp 1435914306
transform 1 0 18720 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_104
timestamp 1435914306
transform 1 0 18720 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_105
timestamp 1435914306
transform 1 0 18720 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_106
timestamp 1435914306
transform 1 0 18720 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_107
timestamp 1435914306
transform 1 0 18720 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_108
timestamp 1435914306
transform 1 0 18720 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_109
timestamp 1435914306
transform 1 0 18720 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_110
timestamp 1435914306
transform 1 0 18720 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_111
timestamp 1435914306
transform 1 0 18720 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_112
timestamp 1435914306
transform 1 0 18720 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_113
timestamp 1435914306
transform 1 0 18720 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_114
timestamp 1435914306
transform 1 0 18720 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_115
timestamp 1435914306
transform 1 0 18720 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_116
timestamp 1435914306
transform 1 0 18720 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_117
timestamp 1435914306
transform 1 0 18720 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_118
timestamp 1435914306
transform 1 0 18720 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_119
timestamp 1435914306
transform 1 0 18720 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_120
timestamp 1435914306
transform 1 0 18720 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_121
timestamp 1435914306
transform 1 0 18720 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_122
timestamp 1435914306
transform 1 0 18720 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_123
timestamp 1435914306
transform 1 0 18720 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_124
timestamp 1435914306
transform 1 0 18720 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_125
timestamp 1435914306
transform 1 0 18720 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_126
timestamp 1435914306
transform 1 0 18720 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_127
timestamp 1435914306
transform 1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_128
timestamp 1435914306
transform -1 0 18720 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_129
timestamp 1435914306
transform -1 0 18720 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_130
timestamp 1435914306
transform -1 0 18720 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_131
timestamp 1435914306
transform -1 0 18720 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_132
timestamp 1435914306
transform -1 0 18720 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_133
timestamp 1435914306
transform -1 0 18720 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_134
timestamp 1435914306
transform -1 0 18720 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_135
timestamp 1435914306
transform -1 0 18720 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_136
timestamp 1435914306
transform -1 0 18720 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_137
timestamp 1435914306
transform -1 0 18720 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_138
timestamp 1435914306
transform -1 0 18720 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_139
timestamp 1435914306
transform -1 0 18720 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_140
timestamp 1435914306
transform -1 0 18720 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_141
timestamp 1435914306
transform -1 0 18720 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_142
timestamp 1435914306
transform -1 0 18720 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_143
timestamp 1435914306
transform -1 0 18720 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_144
timestamp 1435914306
transform -1 0 18720 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_145
timestamp 1435914306
transform -1 0 18720 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_146
timestamp 1435914306
transform -1 0 18720 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_147
timestamp 1435914306
transform -1 0 18720 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_148
timestamp 1435914306
transform -1 0 18720 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_149
timestamp 1435914306
transform -1 0 18720 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_150
timestamp 1435914306
transform -1 0 18720 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_151
timestamp 1435914306
transform -1 0 18720 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_152
timestamp 1435914306
transform -1 0 18720 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_153
timestamp 1435914306
transform -1 0 18720 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_154
timestamp 1435914306
transform -1 0 18720 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_155
timestamp 1435914306
transform -1 0 18720 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_156
timestamp 1435914306
transform -1 0 18720 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_157
timestamp 1435914306
transform -1 0 18720 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_158
timestamp 1435914306
transform -1 0 18720 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_159
timestamp 1435914306
transform -1 0 18720 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_160
timestamp 1435914306
transform -1 0 18720 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_161
timestamp 1435914306
transform -1 0 18720 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_162
timestamp 1435914306
transform -1 0 18720 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_163
timestamp 1435914306
transform -1 0 18720 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_164
timestamp 1435914306
transform -1 0 18720 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_165
timestamp 1435914306
transform -1 0 18720 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_166
timestamp 1435914306
transform -1 0 18720 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_167
timestamp 1435914306
transform -1 0 18720 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_168
timestamp 1435914306
transform -1 0 18720 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_169
timestamp 1435914306
transform -1 0 18720 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_170
timestamp 1435914306
transform -1 0 18720 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_171
timestamp 1435914306
transform -1 0 18720 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_172
timestamp 1435914306
transform -1 0 18720 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_173
timestamp 1435914306
transform -1 0 18720 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_174
timestamp 1435914306
transform -1 0 18720 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_175
timestamp 1435914306
transform -1 0 18720 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_176
timestamp 1435914306
transform -1 0 18720 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_177
timestamp 1435914306
transform -1 0 18720 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_178
timestamp 1435914306
transform -1 0 18720 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_179
timestamp 1435914306
transform -1 0 18720 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_180
timestamp 1435914306
transform -1 0 18720 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_181
timestamp 1435914306
transform -1 0 18720 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_182
timestamp 1435914306
transform -1 0 18720 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_183
timestamp 1435914306
transform -1 0 18720 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_184
timestamp 1435914306
transform -1 0 18720 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_185
timestamp 1435914306
transform -1 0 18720 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_186
timestamp 1435914306
transform -1 0 18720 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_187
timestamp 1435914306
transform -1 0 18720 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_188
timestamp 1435914306
transform -1 0 18720 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_189
timestamp 1435914306
transform -1 0 18720 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_190
timestamp 1435914306
transform -1 0 18720 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_191
timestamp 1435914306
transform -1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_192
timestamp 1435914306
transform 1 0 17472 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_193
timestamp 1435914306
transform 1 0 17472 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_194
timestamp 1435914306
transform 1 0 17472 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_195
timestamp 1435914306
transform 1 0 17472 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_196
timestamp 1435914306
transform 1 0 17472 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_197
timestamp 1435914306
transform 1 0 17472 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_198
timestamp 1435914306
transform 1 0 17472 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_199
timestamp 1435914306
transform 1 0 17472 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_200
timestamp 1435914306
transform 1 0 17472 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_201
timestamp 1435914306
transform 1 0 17472 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_202
timestamp 1435914306
transform 1 0 17472 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_203
timestamp 1435914306
transform 1 0 17472 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_204
timestamp 1435914306
transform 1 0 17472 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_205
timestamp 1435914306
transform 1 0 17472 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_206
timestamp 1435914306
transform 1 0 17472 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_207
timestamp 1435914306
transform 1 0 17472 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_208
timestamp 1435914306
transform 1 0 17472 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_209
timestamp 1435914306
transform 1 0 17472 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_210
timestamp 1435914306
transform 1 0 17472 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_211
timestamp 1435914306
transform 1 0 17472 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_212
timestamp 1435914306
transform 1 0 17472 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_213
timestamp 1435914306
transform 1 0 17472 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_214
timestamp 1435914306
transform 1 0 17472 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_215
timestamp 1435914306
transform 1 0 17472 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_216
timestamp 1435914306
transform 1 0 17472 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_217
timestamp 1435914306
transform 1 0 17472 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_218
timestamp 1435914306
transform 1 0 17472 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_219
timestamp 1435914306
transform 1 0 17472 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_220
timestamp 1435914306
transform 1 0 17472 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_221
timestamp 1435914306
transform 1 0 17472 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_222
timestamp 1435914306
transform 1 0 17472 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_223
timestamp 1435914306
transform 1 0 17472 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_224
timestamp 1435914306
transform 1 0 17472 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_225
timestamp 1435914306
transform 1 0 17472 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_226
timestamp 1435914306
transform 1 0 17472 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_227
timestamp 1435914306
transform 1 0 17472 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_228
timestamp 1435914306
transform 1 0 17472 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_229
timestamp 1435914306
transform 1 0 17472 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_230
timestamp 1435914306
transform 1 0 17472 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_231
timestamp 1435914306
transform 1 0 17472 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_232
timestamp 1435914306
transform 1 0 17472 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_233
timestamp 1435914306
transform 1 0 17472 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_234
timestamp 1435914306
transform 1 0 17472 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_235
timestamp 1435914306
transform 1 0 17472 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_236
timestamp 1435914306
transform 1 0 17472 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_237
timestamp 1435914306
transform 1 0 17472 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_238
timestamp 1435914306
transform 1 0 17472 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_239
timestamp 1435914306
transform 1 0 17472 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_240
timestamp 1435914306
transform 1 0 17472 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_241
timestamp 1435914306
transform 1 0 17472 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_242
timestamp 1435914306
transform 1 0 17472 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_243
timestamp 1435914306
transform 1 0 17472 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_244
timestamp 1435914306
transform 1 0 17472 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_245
timestamp 1435914306
transform 1 0 17472 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_246
timestamp 1435914306
transform 1 0 17472 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_247
timestamp 1435914306
transform 1 0 17472 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_248
timestamp 1435914306
transform 1 0 17472 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_249
timestamp 1435914306
transform 1 0 17472 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_250
timestamp 1435914306
transform 1 0 17472 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_251
timestamp 1435914306
transform 1 0 17472 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_252
timestamp 1435914306
transform 1 0 17472 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_253
timestamp 1435914306
transform 1 0 17472 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_254
timestamp 1435914306
transform 1 0 17472 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_255
timestamp 1435914306
transform 1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_256
timestamp 1435914306
transform -1 0 17472 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_257
timestamp 1435914306
transform -1 0 17472 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_258
timestamp 1435914306
transform -1 0 17472 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_259
timestamp 1435914306
transform -1 0 17472 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_260
timestamp 1435914306
transform -1 0 17472 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_261
timestamp 1435914306
transform -1 0 17472 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_262
timestamp 1435914306
transform -1 0 17472 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_263
timestamp 1435914306
transform -1 0 17472 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_264
timestamp 1435914306
transform -1 0 17472 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_265
timestamp 1435914306
transform -1 0 17472 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_266
timestamp 1435914306
transform -1 0 17472 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_267
timestamp 1435914306
transform -1 0 17472 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_268
timestamp 1435914306
transform -1 0 17472 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_269
timestamp 1435914306
transform -1 0 17472 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_270
timestamp 1435914306
transform -1 0 17472 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_271
timestamp 1435914306
transform -1 0 17472 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_272
timestamp 1435914306
transform -1 0 17472 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_273
timestamp 1435914306
transform -1 0 17472 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_274
timestamp 1435914306
transform -1 0 17472 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_275
timestamp 1435914306
transform -1 0 17472 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_276
timestamp 1435914306
transform -1 0 17472 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_277
timestamp 1435914306
transform -1 0 17472 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_278
timestamp 1435914306
transform -1 0 17472 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_279
timestamp 1435914306
transform -1 0 17472 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_280
timestamp 1435914306
transform -1 0 17472 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_281
timestamp 1435914306
transform -1 0 17472 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_282
timestamp 1435914306
transform -1 0 17472 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_283
timestamp 1435914306
transform -1 0 17472 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_284
timestamp 1435914306
transform -1 0 17472 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_285
timestamp 1435914306
transform -1 0 17472 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_286
timestamp 1435914306
transform -1 0 17472 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_287
timestamp 1435914306
transform -1 0 17472 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_288
timestamp 1435914306
transform -1 0 17472 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_289
timestamp 1435914306
transform -1 0 17472 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_290
timestamp 1435914306
transform -1 0 17472 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_291
timestamp 1435914306
transform -1 0 17472 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_292
timestamp 1435914306
transform -1 0 17472 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_293
timestamp 1435914306
transform -1 0 17472 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_294
timestamp 1435914306
transform -1 0 17472 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_295
timestamp 1435914306
transform -1 0 17472 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_296
timestamp 1435914306
transform -1 0 17472 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_297
timestamp 1435914306
transform -1 0 17472 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_298
timestamp 1435914306
transform -1 0 17472 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_299
timestamp 1435914306
transform -1 0 17472 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_300
timestamp 1435914306
transform -1 0 17472 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_301
timestamp 1435914306
transform -1 0 17472 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_302
timestamp 1435914306
transform -1 0 17472 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_303
timestamp 1435914306
transform -1 0 17472 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_304
timestamp 1435914306
transform -1 0 17472 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_305
timestamp 1435914306
transform -1 0 17472 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_306
timestamp 1435914306
transform -1 0 17472 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_307
timestamp 1435914306
transform -1 0 17472 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_308
timestamp 1435914306
transform -1 0 17472 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_309
timestamp 1435914306
transform -1 0 17472 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_310
timestamp 1435914306
transform -1 0 17472 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_311
timestamp 1435914306
transform -1 0 17472 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_312
timestamp 1435914306
transform -1 0 17472 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_313
timestamp 1435914306
transform -1 0 17472 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_314
timestamp 1435914306
transform -1 0 17472 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_315
timestamp 1435914306
transform -1 0 17472 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_316
timestamp 1435914306
transform -1 0 17472 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_317
timestamp 1435914306
transform -1 0 17472 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_318
timestamp 1435914306
transform -1 0 17472 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_319
timestamp 1435914306
transform -1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_320
timestamp 1435914306
transform 1 0 16224 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_321
timestamp 1435914306
transform 1 0 16224 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_322
timestamp 1435914306
transform 1 0 16224 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_323
timestamp 1435914306
transform 1 0 16224 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_324
timestamp 1435914306
transform 1 0 16224 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_325
timestamp 1435914306
transform 1 0 16224 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_326
timestamp 1435914306
transform 1 0 16224 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_327
timestamp 1435914306
transform 1 0 16224 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_328
timestamp 1435914306
transform 1 0 16224 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_329
timestamp 1435914306
transform 1 0 16224 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_330
timestamp 1435914306
transform 1 0 16224 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_331
timestamp 1435914306
transform 1 0 16224 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_332
timestamp 1435914306
transform 1 0 16224 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_333
timestamp 1435914306
transform 1 0 16224 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_334
timestamp 1435914306
transform 1 0 16224 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_335
timestamp 1435914306
transform 1 0 16224 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_336
timestamp 1435914306
transform 1 0 16224 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_337
timestamp 1435914306
transform 1 0 16224 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_338
timestamp 1435914306
transform 1 0 16224 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_339
timestamp 1435914306
transform 1 0 16224 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_340
timestamp 1435914306
transform 1 0 16224 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_341
timestamp 1435914306
transform 1 0 16224 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_342
timestamp 1435914306
transform 1 0 16224 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_343
timestamp 1435914306
transform 1 0 16224 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_344
timestamp 1435914306
transform 1 0 16224 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_345
timestamp 1435914306
transform 1 0 16224 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_346
timestamp 1435914306
transform 1 0 16224 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_347
timestamp 1435914306
transform 1 0 16224 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_348
timestamp 1435914306
transform 1 0 16224 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_349
timestamp 1435914306
transform 1 0 16224 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_350
timestamp 1435914306
transform 1 0 16224 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_351
timestamp 1435914306
transform 1 0 16224 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_352
timestamp 1435914306
transform 1 0 16224 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_353
timestamp 1435914306
transform 1 0 16224 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_354
timestamp 1435914306
transform 1 0 16224 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_355
timestamp 1435914306
transform 1 0 16224 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_356
timestamp 1435914306
transform 1 0 16224 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_357
timestamp 1435914306
transform 1 0 16224 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_358
timestamp 1435914306
transform 1 0 16224 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_359
timestamp 1435914306
transform 1 0 16224 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_360
timestamp 1435914306
transform 1 0 16224 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_361
timestamp 1435914306
transform 1 0 16224 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_362
timestamp 1435914306
transform 1 0 16224 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_363
timestamp 1435914306
transform 1 0 16224 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_364
timestamp 1435914306
transform 1 0 16224 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_365
timestamp 1435914306
transform 1 0 16224 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_366
timestamp 1435914306
transform 1 0 16224 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_367
timestamp 1435914306
transform 1 0 16224 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_368
timestamp 1435914306
transform 1 0 16224 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_369
timestamp 1435914306
transform 1 0 16224 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_370
timestamp 1435914306
transform 1 0 16224 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_371
timestamp 1435914306
transform 1 0 16224 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_372
timestamp 1435914306
transform 1 0 16224 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_373
timestamp 1435914306
transform 1 0 16224 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_374
timestamp 1435914306
transform 1 0 16224 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_375
timestamp 1435914306
transform 1 0 16224 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_376
timestamp 1435914306
transform 1 0 16224 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_377
timestamp 1435914306
transform 1 0 16224 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_378
timestamp 1435914306
transform 1 0 16224 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_379
timestamp 1435914306
transform 1 0 16224 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_380
timestamp 1435914306
transform 1 0 16224 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_381
timestamp 1435914306
transform 1 0 16224 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_382
timestamp 1435914306
transform 1 0 16224 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_383
timestamp 1435914306
transform 1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_384
timestamp 1435914306
transform -1 0 16224 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_385
timestamp 1435914306
transform -1 0 16224 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_386
timestamp 1435914306
transform -1 0 16224 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_387
timestamp 1435914306
transform -1 0 16224 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_388
timestamp 1435914306
transform -1 0 16224 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_389
timestamp 1435914306
transform -1 0 16224 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_390
timestamp 1435914306
transform -1 0 16224 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_391
timestamp 1435914306
transform -1 0 16224 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_392
timestamp 1435914306
transform -1 0 16224 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_393
timestamp 1435914306
transform -1 0 16224 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_394
timestamp 1435914306
transform -1 0 16224 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_395
timestamp 1435914306
transform -1 0 16224 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_396
timestamp 1435914306
transform -1 0 16224 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_397
timestamp 1435914306
transform -1 0 16224 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_398
timestamp 1435914306
transform -1 0 16224 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_399
timestamp 1435914306
transform -1 0 16224 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_400
timestamp 1435914306
transform -1 0 16224 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_401
timestamp 1435914306
transform -1 0 16224 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_402
timestamp 1435914306
transform -1 0 16224 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_403
timestamp 1435914306
transform -1 0 16224 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_404
timestamp 1435914306
transform -1 0 16224 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_405
timestamp 1435914306
transform -1 0 16224 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_406
timestamp 1435914306
transform -1 0 16224 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_407
timestamp 1435914306
transform -1 0 16224 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_408
timestamp 1435914306
transform -1 0 16224 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_409
timestamp 1435914306
transform -1 0 16224 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_410
timestamp 1435914306
transform -1 0 16224 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_411
timestamp 1435914306
transform -1 0 16224 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_412
timestamp 1435914306
transform -1 0 16224 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_413
timestamp 1435914306
transform -1 0 16224 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_414
timestamp 1435914306
transform -1 0 16224 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_415
timestamp 1435914306
transform -1 0 16224 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_416
timestamp 1435914306
transform -1 0 16224 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_417
timestamp 1435914306
transform -1 0 16224 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_418
timestamp 1435914306
transform -1 0 16224 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_419
timestamp 1435914306
transform -1 0 16224 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_420
timestamp 1435914306
transform -1 0 16224 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_421
timestamp 1435914306
transform -1 0 16224 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_422
timestamp 1435914306
transform -1 0 16224 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_423
timestamp 1435914306
transform -1 0 16224 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_424
timestamp 1435914306
transform -1 0 16224 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_425
timestamp 1435914306
transform -1 0 16224 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_426
timestamp 1435914306
transform -1 0 16224 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_427
timestamp 1435914306
transform -1 0 16224 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_428
timestamp 1435914306
transform -1 0 16224 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_429
timestamp 1435914306
transform -1 0 16224 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_430
timestamp 1435914306
transform -1 0 16224 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_431
timestamp 1435914306
transform -1 0 16224 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_432
timestamp 1435914306
transform -1 0 16224 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_433
timestamp 1435914306
transform -1 0 16224 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_434
timestamp 1435914306
transform -1 0 16224 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_435
timestamp 1435914306
transform -1 0 16224 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_436
timestamp 1435914306
transform -1 0 16224 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_437
timestamp 1435914306
transform -1 0 16224 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_438
timestamp 1435914306
transform -1 0 16224 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_439
timestamp 1435914306
transform -1 0 16224 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_440
timestamp 1435914306
transform -1 0 16224 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_441
timestamp 1435914306
transform -1 0 16224 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_442
timestamp 1435914306
transform -1 0 16224 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_443
timestamp 1435914306
transform -1 0 16224 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_444
timestamp 1435914306
transform -1 0 16224 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_445
timestamp 1435914306
transform -1 0 16224 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_446
timestamp 1435914306
transform -1 0 16224 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_447
timestamp 1435914306
transform -1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_448
timestamp 1435914306
transform 1 0 14976 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_449
timestamp 1435914306
transform 1 0 14976 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_450
timestamp 1435914306
transform 1 0 14976 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_451
timestamp 1435914306
transform 1 0 14976 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_452
timestamp 1435914306
transform 1 0 14976 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_453
timestamp 1435914306
transform 1 0 14976 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_454
timestamp 1435914306
transform 1 0 14976 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_455
timestamp 1435914306
transform 1 0 14976 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_456
timestamp 1435914306
transform 1 0 14976 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_457
timestamp 1435914306
transform 1 0 14976 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_458
timestamp 1435914306
transform 1 0 14976 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_459
timestamp 1435914306
transform 1 0 14976 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_460
timestamp 1435914306
transform 1 0 14976 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_461
timestamp 1435914306
transform 1 0 14976 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_462
timestamp 1435914306
transform 1 0 14976 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_463
timestamp 1435914306
transform 1 0 14976 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_464
timestamp 1435914306
transform 1 0 14976 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_465
timestamp 1435914306
transform 1 0 14976 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_466
timestamp 1435914306
transform 1 0 14976 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_467
timestamp 1435914306
transform 1 0 14976 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_468
timestamp 1435914306
transform 1 0 14976 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_469
timestamp 1435914306
transform 1 0 14976 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_470
timestamp 1435914306
transform 1 0 14976 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_471
timestamp 1435914306
transform 1 0 14976 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_472
timestamp 1435914306
transform 1 0 14976 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_473
timestamp 1435914306
transform 1 0 14976 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_474
timestamp 1435914306
transform 1 0 14976 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_475
timestamp 1435914306
transform 1 0 14976 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_476
timestamp 1435914306
transform 1 0 14976 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_477
timestamp 1435914306
transform 1 0 14976 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_478
timestamp 1435914306
transform 1 0 14976 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_479
timestamp 1435914306
transform 1 0 14976 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_480
timestamp 1435914306
transform 1 0 14976 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_481
timestamp 1435914306
transform 1 0 14976 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_482
timestamp 1435914306
transform 1 0 14976 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_483
timestamp 1435914306
transform 1 0 14976 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_484
timestamp 1435914306
transform 1 0 14976 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_485
timestamp 1435914306
transform 1 0 14976 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_486
timestamp 1435914306
transform 1 0 14976 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_487
timestamp 1435914306
transform 1 0 14976 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_488
timestamp 1435914306
transform 1 0 14976 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_489
timestamp 1435914306
transform 1 0 14976 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_490
timestamp 1435914306
transform 1 0 14976 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_491
timestamp 1435914306
transform 1 0 14976 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_492
timestamp 1435914306
transform 1 0 14976 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_493
timestamp 1435914306
transform 1 0 14976 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_494
timestamp 1435914306
transform 1 0 14976 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_495
timestamp 1435914306
transform 1 0 14976 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_496
timestamp 1435914306
transform 1 0 14976 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_497
timestamp 1435914306
transform 1 0 14976 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_498
timestamp 1435914306
transform 1 0 14976 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_499
timestamp 1435914306
transform 1 0 14976 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_500
timestamp 1435914306
transform 1 0 14976 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_501
timestamp 1435914306
transform 1 0 14976 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_502
timestamp 1435914306
transform 1 0 14976 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_503
timestamp 1435914306
transform 1 0 14976 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_504
timestamp 1435914306
transform 1 0 14976 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_505
timestamp 1435914306
transform 1 0 14976 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_506
timestamp 1435914306
transform 1 0 14976 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_507
timestamp 1435914306
transform 1 0 14976 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_508
timestamp 1435914306
transform 1 0 14976 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_509
timestamp 1435914306
transform 1 0 14976 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_510
timestamp 1435914306
transform 1 0 14976 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_511
timestamp 1435914306
transform 1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_512
timestamp 1435914306
transform -1 0 14976 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_513
timestamp 1435914306
transform -1 0 14976 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_514
timestamp 1435914306
transform -1 0 14976 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_515
timestamp 1435914306
transform -1 0 14976 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_516
timestamp 1435914306
transform -1 0 14976 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_517
timestamp 1435914306
transform -1 0 14976 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_518
timestamp 1435914306
transform -1 0 14976 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_519
timestamp 1435914306
transform -1 0 14976 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_520
timestamp 1435914306
transform -1 0 14976 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_521
timestamp 1435914306
transform -1 0 14976 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_522
timestamp 1435914306
transform -1 0 14976 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_523
timestamp 1435914306
transform -1 0 14976 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_524
timestamp 1435914306
transform -1 0 14976 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_525
timestamp 1435914306
transform -1 0 14976 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_526
timestamp 1435914306
transform -1 0 14976 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_527
timestamp 1435914306
transform -1 0 14976 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_528
timestamp 1435914306
transform -1 0 14976 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_529
timestamp 1435914306
transform -1 0 14976 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_530
timestamp 1435914306
transform -1 0 14976 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_531
timestamp 1435914306
transform -1 0 14976 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_532
timestamp 1435914306
transform -1 0 14976 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_533
timestamp 1435914306
transform -1 0 14976 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_534
timestamp 1435914306
transform -1 0 14976 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_535
timestamp 1435914306
transform -1 0 14976 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_536
timestamp 1435914306
transform -1 0 14976 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_537
timestamp 1435914306
transform -1 0 14976 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_538
timestamp 1435914306
transform -1 0 14976 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_539
timestamp 1435914306
transform -1 0 14976 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_540
timestamp 1435914306
transform -1 0 14976 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_541
timestamp 1435914306
transform -1 0 14976 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_542
timestamp 1435914306
transform -1 0 14976 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_543
timestamp 1435914306
transform -1 0 14976 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_544
timestamp 1435914306
transform -1 0 14976 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_545
timestamp 1435914306
transform -1 0 14976 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_546
timestamp 1435914306
transform -1 0 14976 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_547
timestamp 1435914306
transform -1 0 14976 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_548
timestamp 1435914306
transform -1 0 14976 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_549
timestamp 1435914306
transform -1 0 14976 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_550
timestamp 1435914306
transform -1 0 14976 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_551
timestamp 1435914306
transform -1 0 14976 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_552
timestamp 1435914306
transform -1 0 14976 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_553
timestamp 1435914306
transform -1 0 14976 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_554
timestamp 1435914306
transform -1 0 14976 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_555
timestamp 1435914306
transform -1 0 14976 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_556
timestamp 1435914306
transform -1 0 14976 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_557
timestamp 1435914306
transform -1 0 14976 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_558
timestamp 1435914306
transform -1 0 14976 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_559
timestamp 1435914306
transform -1 0 14976 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_560
timestamp 1435914306
transform -1 0 14976 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_561
timestamp 1435914306
transform -1 0 14976 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_562
timestamp 1435914306
transform -1 0 14976 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_563
timestamp 1435914306
transform -1 0 14976 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_564
timestamp 1435914306
transform -1 0 14976 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_565
timestamp 1435914306
transform -1 0 14976 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_566
timestamp 1435914306
transform -1 0 14976 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_567
timestamp 1435914306
transform -1 0 14976 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_568
timestamp 1435914306
transform -1 0 14976 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_569
timestamp 1435914306
transform -1 0 14976 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_570
timestamp 1435914306
transform -1 0 14976 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_571
timestamp 1435914306
transform -1 0 14976 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_572
timestamp 1435914306
transform -1 0 14976 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_573
timestamp 1435914306
transform -1 0 14976 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_574
timestamp 1435914306
transform -1 0 14976 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_575
timestamp 1435914306
transform -1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_576
timestamp 1435914306
transform 1 0 13728 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_577
timestamp 1435914306
transform 1 0 13728 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_578
timestamp 1435914306
transform 1 0 13728 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_579
timestamp 1435914306
transform 1 0 13728 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_580
timestamp 1435914306
transform 1 0 13728 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_581
timestamp 1435914306
transform 1 0 13728 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_582
timestamp 1435914306
transform 1 0 13728 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_583
timestamp 1435914306
transform 1 0 13728 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_584
timestamp 1435914306
transform 1 0 13728 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_585
timestamp 1435914306
transform 1 0 13728 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_586
timestamp 1435914306
transform 1 0 13728 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_587
timestamp 1435914306
transform 1 0 13728 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_588
timestamp 1435914306
transform 1 0 13728 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_589
timestamp 1435914306
transform 1 0 13728 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_590
timestamp 1435914306
transform 1 0 13728 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_591
timestamp 1435914306
transform 1 0 13728 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_592
timestamp 1435914306
transform 1 0 13728 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_593
timestamp 1435914306
transform 1 0 13728 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_594
timestamp 1435914306
transform 1 0 13728 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_595
timestamp 1435914306
transform 1 0 13728 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_596
timestamp 1435914306
transform 1 0 13728 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_597
timestamp 1435914306
transform 1 0 13728 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_598
timestamp 1435914306
transform 1 0 13728 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_599
timestamp 1435914306
transform 1 0 13728 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_600
timestamp 1435914306
transform 1 0 13728 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_601
timestamp 1435914306
transform 1 0 13728 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_602
timestamp 1435914306
transform 1 0 13728 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_603
timestamp 1435914306
transform 1 0 13728 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_604
timestamp 1435914306
transform 1 0 13728 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_605
timestamp 1435914306
transform 1 0 13728 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_606
timestamp 1435914306
transform 1 0 13728 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_607
timestamp 1435914306
transform 1 0 13728 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_608
timestamp 1435914306
transform 1 0 13728 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_609
timestamp 1435914306
transform 1 0 13728 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_610
timestamp 1435914306
transform 1 0 13728 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_611
timestamp 1435914306
transform 1 0 13728 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_612
timestamp 1435914306
transform 1 0 13728 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_613
timestamp 1435914306
transform 1 0 13728 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_614
timestamp 1435914306
transform 1 0 13728 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_615
timestamp 1435914306
transform 1 0 13728 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_616
timestamp 1435914306
transform 1 0 13728 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_617
timestamp 1435914306
transform 1 0 13728 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_618
timestamp 1435914306
transform 1 0 13728 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_619
timestamp 1435914306
transform 1 0 13728 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_620
timestamp 1435914306
transform 1 0 13728 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_621
timestamp 1435914306
transform 1 0 13728 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_622
timestamp 1435914306
transform 1 0 13728 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_623
timestamp 1435914306
transform 1 0 13728 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_624
timestamp 1435914306
transform 1 0 13728 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_625
timestamp 1435914306
transform 1 0 13728 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_626
timestamp 1435914306
transform 1 0 13728 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_627
timestamp 1435914306
transform 1 0 13728 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_628
timestamp 1435914306
transform 1 0 13728 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_629
timestamp 1435914306
transform 1 0 13728 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_630
timestamp 1435914306
transform 1 0 13728 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_631
timestamp 1435914306
transform 1 0 13728 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_632
timestamp 1435914306
transform 1 0 13728 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_633
timestamp 1435914306
transform 1 0 13728 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_634
timestamp 1435914306
transform 1 0 13728 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_635
timestamp 1435914306
transform 1 0 13728 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_636
timestamp 1435914306
transform 1 0 13728 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_637
timestamp 1435914306
transform 1 0 13728 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_638
timestamp 1435914306
transform 1 0 13728 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_639
timestamp 1435914306
transform 1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_640
timestamp 1435914306
transform -1 0 13728 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_641
timestamp 1435914306
transform -1 0 13728 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_642
timestamp 1435914306
transform -1 0 13728 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_643
timestamp 1435914306
transform -1 0 13728 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_644
timestamp 1435914306
transform -1 0 13728 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_645
timestamp 1435914306
transform -1 0 13728 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_646
timestamp 1435914306
transform -1 0 13728 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_647
timestamp 1435914306
transform -1 0 13728 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_648
timestamp 1435914306
transform -1 0 13728 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_649
timestamp 1435914306
transform -1 0 13728 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_650
timestamp 1435914306
transform -1 0 13728 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_651
timestamp 1435914306
transform -1 0 13728 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_652
timestamp 1435914306
transform -1 0 13728 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_653
timestamp 1435914306
transform -1 0 13728 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_654
timestamp 1435914306
transform -1 0 13728 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_655
timestamp 1435914306
transform -1 0 13728 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_656
timestamp 1435914306
transform -1 0 13728 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_657
timestamp 1435914306
transform -1 0 13728 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_658
timestamp 1435914306
transform -1 0 13728 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_659
timestamp 1435914306
transform -1 0 13728 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_660
timestamp 1435914306
transform -1 0 13728 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_661
timestamp 1435914306
transform -1 0 13728 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_662
timestamp 1435914306
transform -1 0 13728 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_663
timestamp 1435914306
transform -1 0 13728 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_664
timestamp 1435914306
transform -1 0 13728 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_665
timestamp 1435914306
transform -1 0 13728 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_666
timestamp 1435914306
transform -1 0 13728 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_667
timestamp 1435914306
transform -1 0 13728 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_668
timestamp 1435914306
transform -1 0 13728 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_669
timestamp 1435914306
transform -1 0 13728 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_670
timestamp 1435914306
transform -1 0 13728 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_671
timestamp 1435914306
transform -1 0 13728 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_672
timestamp 1435914306
transform -1 0 13728 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_673
timestamp 1435914306
transform -1 0 13728 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_674
timestamp 1435914306
transform -1 0 13728 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_675
timestamp 1435914306
transform -1 0 13728 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_676
timestamp 1435914306
transform -1 0 13728 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_677
timestamp 1435914306
transform -1 0 13728 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_678
timestamp 1435914306
transform -1 0 13728 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_679
timestamp 1435914306
transform -1 0 13728 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_680
timestamp 1435914306
transform -1 0 13728 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_681
timestamp 1435914306
transform -1 0 13728 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_682
timestamp 1435914306
transform -1 0 13728 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_683
timestamp 1435914306
transform -1 0 13728 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_684
timestamp 1435914306
transform -1 0 13728 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_685
timestamp 1435914306
transform -1 0 13728 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_686
timestamp 1435914306
transform -1 0 13728 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_687
timestamp 1435914306
transform -1 0 13728 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_688
timestamp 1435914306
transform -1 0 13728 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_689
timestamp 1435914306
transform -1 0 13728 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_690
timestamp 1435914306
transform -1 0 13728 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_691
timestamp 1435914306
transform -1 0 13728 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_692
timestamp 1435914306
transform -1 0 13728 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_693
timestamp 1435914306
transform -1 0 13728 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_694
timestamp 1435914306
transform -1 0 13728 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_695
timestamp 1435914306
transform -1 0 13728 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_696
timestamp 1435914306
transform -1 0 13728 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_697
timestamp 1435914306
transform -1 0 13728 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_698
timestamp 1435914306
transform -1 0 13728 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_699
timestamp 1435914306
transform -1 0 13728 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_700
timestamp 1435914306
transform -1 0 13728 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_701
timestamp 1435914306
transform -1 0 13728 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_702
timestamp 1435914306
transform -1 0 13728 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_703
timestamp 1435914306
transform -1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_704
timestamp 1435914306
transform 1 0 12480 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_705
timestamp 1435914306
transform 1 0 12480 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_706
timestamp 1435914306
transform 1 0 12480 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_707
timestamp 1435914306
transform 1 0 12480 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_708
timestamp 1435914306
transform 1 0 12480 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_709
timestamp 1435914306
transform 1 0 12480 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_710
timestamp 1435914306
transform 1 0 12480 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_711
timestamp 1435914306
transform 1 0 12480 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_712
timestamp 1435914306
transform 1 0 12480 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_713
timestamp 1435914306
transform 1 0 12480 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_714
timestamp 1435914306
transform 1 0 12480 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_715
timestamp 1435914306
transform 1 0 12480 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_716
timestamp 1435914306
transform 1 0 12480 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_717
timestamp 1435914306
transform 1 0 12480 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_718
timestamp 1435914306
transform 1 0 12480 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_719
timestamp 1435914306
transform 1 0 12480 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_720
timestamp 1435914306
transform 1 0 12480 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_721
timestamp 1435914306
transform 1 0 12480 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_722
timestamp 1435914306
transform 1 0 12480 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_723
timestamp 1435914306
transform 1 0 12480 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_724
timestamp 1435914306
transform 1 0 12480 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_725
timestamp 1435914306
transform 1 0 12480 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_726
timestamp 1435914306
transform 1 0 12480 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_727
timestamp 1435914306
transform 1 0 12480 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_728
timestamp 1435914306
transform 1 0 12480 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_729
timestamp 1435914306
transform 1 0 12480 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_730
timestamp 1435914306
transform 1 0 12480 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_731
timestamp 1435914306
transform 1 0 12480 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_732
timestamp 1435914306
transform 1 0 12480 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_733
timestamp 1435914306
transform 1 0 12480 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_734
timestamp 1435914306
transform 1 0 12480 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_735
timestamp 1435914306
transform 1 0 12480 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_736
timestamp 1435914306
transform 1 0 12480 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_737
timestamp 1435914306
transform 1 0 12480 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_738
timestamp 1435914306
transform 1 0 12480 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_739
timestamp 1435914306
transform 1 0 12480 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_740
timestamp 1435914306
transform 1 0 12480 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_741
timestamp 1435914306
transform 1 0 12480 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_742
timestamp 1435914306
transform 1 0 12480 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_743
timestamp 1435914306
transform 1 0 12480 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_744
timestamp 1435914306
transform 1 0 12480 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_745
timestamp 1435914306
transform 1 0 12480 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_746
timestamp 1435914306
transform 1 0 12480 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_747
timestamp 1435914306
transform 1 0 12480 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_748
timestamp 1435914306
transform 1 0 12480 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_749
timestamp 1435914306
transform 1 0 12480 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_750
timestamp 1435914306
transform 1 0 12480 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_751
timestamp 1435914306
transform 1 0 12480 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_752
timestamp 1435914306
transform 1 0 12480 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_753
timestamp 1435914306
transform 1 0 12480 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_754
timestamp 1435914306
transform 1 0 12480 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_755
timestamp 1435914306
transform 1 0 12480 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_756
timestamp 1435914306
transform 1 0 12480 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_757
timestamp 1435914306
transform 1 0 12480 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_758
timestamp 1435914306
transform 1 0 12480 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_759
timestamp 1435914306
transform 1 0 12480 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_760
timestamp 1435914306
transform 1 0 12480 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_761
timestamp 1435914306
transform 1 0 12480 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_762
timestamp 1435914306
transform 1 0 12480 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_763
timestamp 1435914306
transform 1 0 12480 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_764
timestamp 1435914306
transform 1 0 12480 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_765
timestamp 1435914306
transform 1 0 12480 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_766
timestamp 1435914306
transform 1 0 12480 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_767
timestamp 1435914306
transform 1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_768
timestamp 1435914306
transform -1 0 12480 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_769
timestamp 1435914306
transform -1 0 12480 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_770
timestamp 1435914306
transform -1 0 12480 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_771
timestamp 1435914306
transform -1 0 12480 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_772
timestamp 1435914306
transform -1 0 12480 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_773
timestamp 1435914306
transform -1 0 12480 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_774
timestamp 1435914306
transform -1 0 12480 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_775
timestamp 1435914306
transform -1 0 12480 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_776
timestamp 1435914306
transform -1 0 12480 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_777
timestamp 1435914306
transform -1 0 12480 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_778
timestamp 1435914306
transform -1 0 12480 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_779
timestamp 1435914306
transform -1 0 12480 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_780
timestamp 1435914306
transform -1 0 12480 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_781
timestamp 1435914306
transform -1 0 12480 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_782
timestamp 1435914306
transform -1 0 12480 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_783
timestamp 1435914306
transform -1 0 12480 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_784
timestamp 1435914306
transform -1 0 12480 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_785
timestamp 1435914306
transform -1 0 12480 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_786
timestamp 1435914306
transform -1 0 12480 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_787
timestamp 1435914306
transform -1 0 12480 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_788
timestamp 1435914306
transform -1 0 12480 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_789
timestamp 1435914306
transform -1 0 12480 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_790
timestamp 1435914306
transform -1 0 12480 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_791
timestamp 1435914306
transform -1 0 12480 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_792
timestamp 1435914306
transform -1 0 12480 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_793
timestamp 1435914306
transform -1 0 12480 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_794
timestamp 1435914306
transform -1 0 12480 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_795
timestamp 1435914306
transform -1 0 12480 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_796
timestamp 1435914306
transform -1 0 12480 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_797
timestamp 1435914306
transform -1 0 12480 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_798
timestamp 1435914306
transform -1 0 12480 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_799
timestamp 1435914306
transform -1 0 12480 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_800
timestamp 1435914306
transform -1 0 12480 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_801
timestamp 1435914306
transform -1 0 12480 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_802
timestamp 1435914306
transform -1 0 12480 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_803
timestamp 1435914306
transform -1 0 12480 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_804
timestamp 1435914306
transform -1 0 12480 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_805
timestamp 1435914306
transform -1 0 12480 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_806
timestamp 1435914306
transform -1 0 12480 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_807
timestamp 1435914306
transform -1 0 12480 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_808
timestamp 1435914306
transform -1 0 12480 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_809
timestamp 1435914306
transform -1 0 12480 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_810
timestamp 1435914306
transform -1 0 12480 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_811
timestamp 1435914306
transform -1 0 12480 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_812
timestamp 1435914306
transform -1 0 12480 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_813
timestamp 1435914306
transform -1 0 12480 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_814
timestamp 1435914306
transform -1 0 12480 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_815
timestamp 1435914306
transform -1 0 12480 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_816
timestamp 1435914306
transform -1 0 12480 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_817
timestamp 1435914306
transform -1 0 12480 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_818
timestamp 1435914306
transform -1 0 12480 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_819
timestamp 1435914306
transform -1 0 12480 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_820
timestamp 1435914306
transform -1 0 12480 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_821
timestamp 1435914306
transform -1 0 12480 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_822
timestamp 1435914306
transform -1 0 12480 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_823
timestamp 1435914306
transform -1 0 12480 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_824
timestamp 1435914306
transform -1 0 12480 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_825
timestamp 1435914306
transform -1 0 12480 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_826
timestamp 1435914306
transform -1 0 12480 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_827
timestamp 1435914306
transform -1 0 12480 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_828
timestamp 1435914306
transform -1 0 12480 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_829
timestamp 1435914306
transform -1 0 12480 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_830
timestamp 1435914306
transform -1 0 12480 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_831
timestamp 1435914306
transform -1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_832
timestamp 1435914306
transform 1 0 11232 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_833
timestamp 1435914306
transform 1 0 11232 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_834
timestamp 1435914306
transform 1 0 11232 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_835
timestamp 1435914306
transform 1 0 11232 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_836
timestamp 1435914306
transform 1 0 11232 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_837
timestamp 1435914306
transform 1 0 11232 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_838
timestamp 1435914306
transform 1 0 11232 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_839
timestamp 1435914306
transform 1 0 11232 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_840
timestamp 1435914306
transform 1 0 11232 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_841
timestamp 1435914306
transform 1 0 11232 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_842
timestamp 1435914306
transform 1 0 11232 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_843
timestamp 1435914306
transform 1 0 11232 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_844
timestamp 1435914306
transform 1 0 11232 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_845
timestamp 1435914306
transform 1 0 11232 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_846
timestamp 1435914306
transform 1 0 11232 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_847
timestamp 1435914306
transform 1 0 11232 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_848
timestamp 1435914306
transform 1 0 11232 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_849
timestamp 1435914306
transform 1 0 11232 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_850
timestamp 1435914306
transform 1 0 11232 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_851
timestamp 1435914306
transform 1 0 11232 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_852
timestamp 1435914306
transform 1 0 11232 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_853
timestamp 1435914306
transform 1 0 11232 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_854
timestamp 1435914306
transform 1 0 11232 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_855
timestamp 1435914306
transform 1 0 11232 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_856
timestamp 1435914306
transform 1 0 11232 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_857
timestamp 1435914306
transform 1 0 11232 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_858
timestamp 1435914306
transform 1 0 11232 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_859
timestamp 1435914306
transform 1 0 11232 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_860
timestamp 1435914306
transform 1 0 11232 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_861
timestamp 1435914306
transform 1 0 11232 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_862
timestamp 1435914306
transform 1 0 11232 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_863
timestamp 1435914306
transform 1 0 11232 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_864
timestamp 1435914306
transform 1 0 11232 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_865
timestamp 1435914306
transform 1 0 11232 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_866
timestamp 1435914306
transform 1 0 11232 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_867
timestamp 1435914306
transform 1 0 11232 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_868
timestamp 1435914306
transform 1 0 11232 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_869
timestamp 1435914306
transform 1 0 11232 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_870
timestamp 1435914306
transform 1 0 11232 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_871
timestamp 1435914306
transform 1 0 11232 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_872
timestamp 1435914306
transform 1 0 11232 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_873
timestamp 1435914306
transform 1 0 11232 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_874
timestamp 1435914306
transform 1 0 11232 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_875
timestamp 1435914306
transform 1 0 11232 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_876
timestamp 1435914306
transform 1 0 11232 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_877
timestamp 1435914306
transform 1 0 11232 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_878
timestamp 1435914306
transform 1 0 11232 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_879
timestamp 1435914306
transform 1 0 11232 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_880
timestamp 1435914306
transform 1 0 11232 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_881
timestamp 1435914306
transform 1 0 11232 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_882
timestamp 1435914306
transform 1 0 11232 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_883
timestamp 1435914306
transform 1 0 11232 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_884
timestamp 1435914306
transform 1 0 11232 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_885
timestamp 1435914306
transform 1 0 11232 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_886
timestamp 1435914306
transform 1 0 11232 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_887
timestamp 1435914306
transform 1 0 11232 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_888
timestamp 1435914306
transform 1 0 11232 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_889
timestamp 1435914306
transform 1 0 11232 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_890
timestamp 1435914306
transform 1 0 11232 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_891
timestamp 1435914306
transform 1 0 11232 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_892
timestamp 1435914306
transform 1 0 11232 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_893
timestamp 1435914306
transform 1 0 11232 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_894
timestamp 1435914306
transform 1 0 11232 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_895
timestamp 1435914306
transform 1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_896
timestamp 1435914306
transform -1 0 11232 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_897
timestamp 1435914306
transform -1 0 11232 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_898
timestamp 1435914306
transform -1 0 11232 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_899
timestamp 1435914306
transform -1 0 11232 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_900
timestamp 1435914306
transform -1 0 11232 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_901
timestamp 1435914306
transform -1 0 11232 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_902
timestamp 1435914306
transform -1 0 11232 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_903
timestamp 1435914306
transform -1 0 11232 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_904
timestamp 1435914306
transform -1 0 11232 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_905
timestamp 1435914306
transform -1 0 11232 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_906
timestamp 1435914306
transform -1 0 11232 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_907
timestamp 1435914306
transform -1 0 11232 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_908
timestamp 1435914306
transform -1 0 11232 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_909
timestamp 1435914306
transform -1 0 11232 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_910
timestamp 1435914306
transform -1 0 11232 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_911
timestamp 1435914306
transform -1 0 11232 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_912
timestamp 1435914306
transform -1 0 11232 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_913
timestamp 1435914306
transform -1 0 11232 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_914
timestamp 1435914306
transform -1 0 11232 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_915
timestamp 1435914306
transform -1 0 11232 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_916
timestamp 1435914306
transform -1 0 11232 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_917
timestamp 1435914306
transform -1 0 11232 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_918
timestamp 1435914306
transform -1 0 11232 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_919
timestamp 1435914306
transform -1 0 11232 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_920
timestamp 1435914306
transform -1 0 11232 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_921
timestamp 1435914306
transform -1 0 11232 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_922
timestamp 1435914306
transform -1 0 11232 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_923
timestamp 1435914306
transform -1 0 11232 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_924
timestamp 1435914306
transform -1 0 11232 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_925
timestamp 1435914306
transform -1 0 11232 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_926
timestamp 1435914306
transform -1 0 11232 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_927
timestamp 1435914306
transform -1 0 11232 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_928
timestamp 1435914306
transform -1 0 11232 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_929
timestamp 1435914306
transform -1 0 11232 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_930
timestamp 1435914306
transform -1 0 11232 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_931
timestamp 1435914306
transform -1 0 11232 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_932
timestamp 1435914306
transform -1 0 11232 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_933
timestamp 1435914306
transform -1 0 11232 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_934
timestamp 1435914306
transform -1 0 11232 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_935
timestamp 1435914306
transform -1 0 11232 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_936
timestamp 1435914306
transform -1 0 11232 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_937
timestamp 1435914306
transform -1 0 11232 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_938
timestamp 1435914306
transform -1 0 11232 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_939
timestamp 1435914306
transform -1 0 11232 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_940
timestamp 1435914306
transform -1 0 11232 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_941
timestamp 1435914306
transform -1 0 11232 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_942
timestamp 1435914306
transform -1 0 11232 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_943
timestamp 1435914306
transform -1 0 11232 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_944
timestamp 1435914306
transform -1 0 11232 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_945
timestamp 1435914306
transform -1 0 11232 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_946
timestamp 1435914306
transform -1 0 11232 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_947
timestamp 1435914306
transform -1 0 11232 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_948
timestamp 1435914306
transform -1 0 11232 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_949
timestamp 1435914306
transform -1 0 11232 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_950
timestamp 1435914306
transform -1 0 11232 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_951
timestamp 1435914306
transform -1 0 11232 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_952
timestamp 1435914306
transform -1 0 11232 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_953
timestamp 1435914306
transform -1 0 11232 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_954
timestamp 1435914306
transform -1 0 11232 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_955
timestamp 1435914306
transform -1 0 11232 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_956
timestamp 1435914306
transform -1 0 11232 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_957
timestamp 1435914306
transform -1 0 11232 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_958
timestamp 1435914306
transform -1 0 11232 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_959
timestamp 1435914306
transform -1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_960
timestamp 1435914306
transform 1 0 9984 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_961
timestamp 1435914306
transform 1 0 9984 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_962
timestamp 1435914306
transform 1 0 9984 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_963
timestamp 1435914306
transform 1 0 9984 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_964
timestamp 1435914306
transform 1 0 9984 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_965
timestamp 1435914306
transform 1 0 9984 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_966
timestamp 1435914306
transform 1 0 9984 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_967
timestamp 1435914306
transform 1 0 9984 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_968
timestamp 1435914306
transform 1 0 9984 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_969
timestamp 1435914306
transform 1 0 9984 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_970
timestamp 1435914306
transform 1 0 9984 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_971
timestamp 1435914306
transform 1 0 9984 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_972
timestamp 1435914306
transform 1 0 9984 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_973
timestamp 1435914306
transform 1 0 9984 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_974
timestamp 1435914306
transform 1 0 9984 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_975
timestamp 1435914306
transform 1 0 9984 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_976
timestamp 1435914306
transform 1 0 9984 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_977
timestamp 1435914306
transform 1 0 9984 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_978
timestamp 1435914306
transform 1 0 9984 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_979
timestamp 1435914306
transform 1 0 9984 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_980
timestamp 1435914306
transform 1 0 9984 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_981
timestamp 1435914306
transform 1 0 9984 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_982
timestamp 1435914306
transform 1 0 9984 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_983
timestamp 1435914306
transform 1 0 9984 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_984
timestamp 1435914306
transform 1 0 9984 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_985
timestamp 1435914306
transform 1 0 9984 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_986
timestamp 1435914306
transform 1 0 9984 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_987
timestamp 1435914306
transform 1 0 9984 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_988
timestamp 1435914306
transform 1 0 9984 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_989
timestamp 1435914306
transform 1 0 9984 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_990
timestamp 1435914306
transform 1 0 9984 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_991
timestamp 1435914306
transform 1 0 9984 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_992
timestamp 1435914306
transform 1 0 9984 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_993
timestamp 1435914306
transform 1 0 9984 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_994
timestamp 1435914306
transform 1 0 9984 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_995
timestamp 1435914306
transform 1 0 9984 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_996
timestamp 1435914306
transform 1 0 9984 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_997
timestamp 1435914306
transform 1 0 9984 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_998
timestamp 1435914306
transform 1 0 9984 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_999
timestamp 1435914306
transform 1 0 9984 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1000
timestamp 1435914306
transform 1 0 9984 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1001
timestamp 1435914306
transform 1 0 9984 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1002
timestamp 1435914306
transform 1 0 9984 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1003
timestamp 1435914306
transform 1 0 9984 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1004
timestamp 1435914306
transform 1 0 9984 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1005
timestamp 1435914306
transform 1 0 9984 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1006
timestamp 1435914306
transform 1 0 9984 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1007
timestamp 1435914306
transform 1 0 9984 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1008
timestamp 1435914306
transform 1 0 9984 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1009
timestamp 1435914306
transform 1 0 9984 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1010
timestamp 1435914306
transform 1 0 9984 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1011
timestamp 1435914306
transform 1 0 9984 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1012
timestamp 1435914306
transform 1 0 9984 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1013
timestamp 1435914306
transform 1 0 9984 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1014
timestamp 1435914306
transform 1 0 9984 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1015
timestamp 1435914306
transform 1 0 9984 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1016
timestamp 1435914306
transform 1 0 9984 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1017
timestamp 1435914306
transform 1 0 9984 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1018
timestamp 1435914306
transform 1 0 9984 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1019
timestamp 1435914306
transform 1 0 9984 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1020
timestamp 1435914306
transform 1 0 9984 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1021
timestamp 1435914306
transform 1 0 9984 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1022
timestamp 1435914306
transform 1 0 9984 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1023
timestamp 1435914306
transform 1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1024
timestamp 1435914306
transform -1 0 9984 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1025
timestamp 1435914306
transform -1 0 9984 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1026
timestamp 1435914306
transform -1 0 9984 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1027
timestamp 1435914306
transform -1 0 9984 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1028
timestamp 1435914306
transform -1 0 9984 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1029
timestamp 1435914306
transform -1 0 9984 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1030
timestamp 1435914306
transform -1 0 9984 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1031
timestamp 1435914306
transform -1 0 9984 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1032
timestamp 1435914306
transform -1 0 9984 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1033
timestamp 1435914306
transform -1 0 9984 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1034
timestamp 1435914306
transform -1 0 9984 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1035
timestamp 1435914306
transform -1 0 9984 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1036
timestamp 1435914306
transform -1 0 9984 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1037
timestamp 1435914306
transform -1 0 9984 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1038
timestamp 1435914306
transform -1 0 9984 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1039
timestamp 1435914306
transform -1 0 9984 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1040
timestamp 1435914306
transform -1 0 9984 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1041
timestamp 1435914306
transform -1 0 9984 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1042
timestamp 1435914306
transform -1 0 9984 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1043
timestamp 1435914306
transform -1 0 9984 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1044
timestamp 1435914306
transform -1 0 9984 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1045
timestamp 1435914306
transform -1 0 9984 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1046
timestamp 1435914306
transform -1 0 9984 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1047
timestamp 1435914306
transform -1 0 9984 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1048
timestamp 1435914306
transform -1 0 9984 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1049
timestamp 1435914306
transform -1 0 9984 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1050
timestamp 1435914306
transform -1 0 9984 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1051
timestamp 1435914306
transform -1 0 9984 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1052
timestamp 1435914306
transform -1 0 9984 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1053
timestamp 1435914306
transform -1 0 9984 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1054
timestamp 1435914306
transform -1 0 9984 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1055
timestamp 1435914306
transform -1 0 9984 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1056
timestamp 1435914306
transform -1 0 9984 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1057
timestamp 1435914306
transform -1 0 9984 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1058
timestamp 1435914306
transform -1 0 9984 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1059
timestamp 1435914306
transform -1 0 9984 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1060
timestamp 1435914306
transform -1 0 9984 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1061
timestamp 1435914306
transform -1 0 9984 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1062
timestamp 1435914306
transform -1 0 9984 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1063
timestamp 1435914306
transform -1 0 9984 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1064
timestamp 1435914306
transform -1 0 9984 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1065
timestamp 1435914306
transform -1 0 9984 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1066
timestamp 1435914306
transform -1 0 9984 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1067
timestamp 1435914306
transform -1 0 9984 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1068
timestamp 1435914306
transform -1 0 9984 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1069
timestamp 1435914306
transform -1 0 9984 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1070
timestamp 1435914306
transform -1 0 9984 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1071
timestamp 1435914306
transform -1 0 9984 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1072
timestamp 1435914306
transform -1 0 9984 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1073
timestamp 1435914306
transform -1 0 9984 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1074
timestamp 1435914306
transform -1 0 9984 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1075
timestamp 1435914306
transform -1 0 9984 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1076
timestamp 1435914306
transform -1 0 9984 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1077
timestamp 1435914306
transform -1 0 9984 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1078
timestamp 1435914306
transform -1 0 9984 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1079
timestamp 1435914306
transform -1 0 9984 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1080
timestamp 1435914306
transform -1 0 9984 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1081
timestamp 1435914306
transform -1 0 9984 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1082
timestamp 1435914306
transform -1 0 9984 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1083
timestamp 1435914306
transform -1 0 9984 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1084
timestamp 1435914306
transform -1 0 9984 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1085
timestamp 1435914306
transform -1 0 9984 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1086
timestamp 1435914306
transform -1 0 9984 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1087
timestamp 1435914306
transform -1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1088
timestamp 1435914306
transform 1 0 8736 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1089
timestamp 1435914306
transform 1 0 8736 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1090
timestamp 1435914306
transform 1 0 8736 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1091
timestamp 1435914306
transform 1 0 8736 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1092
timestamp 1435914306
transform 1 0 8736 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1093
timestamp 1435914306
transform 1 0 8736 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1094
timestamp 1435914306
transform 1 0 8736 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1095
timestamp 1435914306
transform 1 0 8736 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1096
timestamp 1435914306
transform 1 0 8736 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1097
timestamp 1435914306
transform 1 0 8736 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1098
timestamp 1435914306
transform 1 0 8736 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1099
timestamp 1435914306
transform 1 0 8736 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1100
timestamp 1435914306
transform 1 0 8736 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1101
timestamp 1435914306
transform 1 0 8736 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1102
timestamp 1435914306
transform 1 0 8736 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1103
timestamp 1435914306
transform 1 0 8736 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1104
timestamp 1435914306
transform 1 0 8736 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1105
timestamp 1435914306
transform 1 0 8736 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1106
timestamp 1435914306
transform 1 0 8736 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1107
timestamp 1435914306
transform 1 0 8736 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1108
timestamp 1435914306
transform 1 0 8736 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1109
timestamp 1435914306
transform 1 0 8736 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1110
timestamp 1435914306
transform 1 0 8736 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1111
timestamp 1435914306
transform 1 0 8736 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1112
timestamp 1435914306
transform 1 0 8736 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1113
timestamp 1435914306
transform 1 0 8736 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1114
timestamp 1435914306
transform 1 0 8736 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1115
timestamp 1435914306
transform 1 0 8736 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1116
timestamp 1435914306
transform 1 0 8736 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1117
timestamp 1435914306
transform 1 0 8736 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1118
timestamp 1435914306
transform 1 0 8736 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1119
timestamp 1435914306
transform 1 0 8736 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1120
timestamp 1435914306
transform 1 0 8736 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1121
timestamp 1435914306
transform 1 0 8736 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1122
timestamp 1435914306
transform 1 0 8736 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1123
timestamp 1435914306
transform 1 0 8736 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1124
timestamp 1435914306
transform 1 0 8736 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1125
timestamp 1435914306
transform 1 0 8736 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1126
timestamp 1435914306
transform 1 0 8736 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1127
timestamp 1435914306
transform 1 0 8736 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1128
timestamp 1435914306
transform 1 0 8736 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1129
timestamp 1435914306
transform 1 0 8736 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1130
timestamp 1435914306
transform 1 0 8736 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1131
timestamp 1435914306
transform 1 0 8736 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1132
timestamp 1435914306
transform 1 0 8736 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1133
timestamp 1435914306
transform 1 0 8736 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1134
timestamp 1435914306
transform 1 0 8736 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1135
timestamp 1435914306
transform 1 0 8736 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1136
timestamp 1435914306
transform 1 0 8736 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1137
timestamp 1435914306
transform 1 0 8736 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1138
timestamp 1435914306
transform 1 0 8736 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1139
timestamp 1435914306
transform 1 0 8736 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1140
timestamp 1435914306
transform 1 0 8736 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1141
timestamp 1435914306
transform 1 0 8736 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1142
timestamp 1435914306
transform 1 0 8736 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1143
timestamp 1435914306
transform 1 0 8736 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1144
timestamp 1435914306
transform 1 0 8736 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1145
timestamp 1435914306
transform 1 0 8736 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1146
timestamp 1435914306
transform 1 0 8736 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1147
timestamp 1435914306
transform 1 0 8736 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1148
timestamp 1435914306
transform 1 0 8736 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1149
timestamp 1435914306
transform 1 0 8736 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1150
timestamp 1435914306
transform 1 0 8736 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1151
timestamp 1435914306
transform 1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1152
timestamp 1435914306
transform -1 0 8736 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1153
timestamp 1435914306
transform -1 0 8736 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1154
timestamp 1435914306
transform -1 0 8736 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1155
timestamp 1435914306
transform -1 0 8736 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1156
timestamp 1435914306
transform -1 0 8736 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1157
timestamp 1435914306
transform -1 0 8736 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1158
timestamp 1435914306
transform -1 0 8736 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1159
timestamp 1435914306
transform -1 0 8736 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1160
timestamp 1435914306
transform -1 0 8736 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1161
timestamp 1435914306
transform -1 0 8736 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1162
timestamp 1435914306
transform -1 0 8736 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1163
timestamp 1435914306
transform -1 0 8736 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1164
timestamp 1435914306
transform -1 0 8736 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1165
timestamp 1435914306
transform -1 0 8736 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1166
timestamp 1435914306
transform -1 0 8736 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1167
timestamp 1435914306
transform -1 0 8736 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1168
timestamp 1435914306
transform -1 0 8736 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1169
timestamp 1435914306
transform -1 0 8736 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1170
timestamp 1435914306
transform -1 0 8736 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1171
timestamp 1435914306
transform -1 0 8736 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1172
timestamp 1435914306
transform -1 0 8736 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1173
timestamp 1435914306
transform -1 0 8736 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1174
timestamp 1435914306
transform -1 0 8736 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1175
timestamp 1435914306
transform -1 0 8736 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1176
timestamp 1435914306
transform -1 0 8736 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1177
timestamp 1435914306
transform -1 0 8736 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1178
timestamp 1435914306
transform -1 0 8736 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1179
timestamp 1435914306
transform -1 0 8736 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1180
timestamp 1435914306
transform -1 0 8736 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1181
timestamp 1435914306
transform -1 0 8736 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1182
timestamp 1435914306
transform -1 0 8736 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1183
timestamp 1435914306
transform -1 0 8736 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1184
timestamp 1435914306
transform -1 0 8736 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1185
timestamp 1435914306
transform -1 0 8736 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1186
timestamp 1435914306
transform -1 0 8736 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1187
timestamp 1435914306
transform -1 0 8736 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1188
timestamp 1435914306
transform -1 0 8736 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1189
timestamp 1435914306
transform -1 0 8736 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1190
timestamp 1435914306
transform -1 0 8736 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1191
timestamp 1435914306
transform -1 0 8736 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1192
timestamp 1435914306
transform -1 0 8736 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1193
timestamp 1435914306
transform -1 0 8736 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1194
timestamp 1435914306
transform -1 0 8736 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1195
timestamp 1435914306
transform -1 0 8736 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1196
timestamp 1435914306
transform -1 0 8736 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1197
timestamp 1435914306
transform -1 0 8736 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1198
timestamp 1435914306
transform -1 0 8736 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1199
timestamp 1435914306
transform -1 0 8736 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1200
timestamp 1435914306
transform -1 0 8736 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1201
timestamp 1435914306
transform -1 0 8736 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1202
timestamp 1435914306
transform -1 0 8736 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1203
timestamp 1435914306
transform -1 0 8736 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1204
timestamp 1435914306
transform -1 0 8736 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1205
timestamp 1435914306
transform -1 0 8736 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1206
timestamp 1435914306
transform -1 0 8736 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1207
timestamp 1435914306
transform -1 0 8736 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1208
timestamp 1435914306
transform -1 0 8736 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1209
timestamp 1435914306
transform -1 0 8736 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1210
timestamp 1435914306
transform -1 0 8736 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1211
timestamp 1435914306
transform -1 0 8736 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1212
timestamp 1435914306
transform -1 0 8736 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1213
timestamp 1435914306
transform -1 0 8736 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1214
timestamp 1435914306
transform -1 0 8736 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1215
timestamp 1435914306
transform -1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1216
timestamp 1435914306
transform 1 0 7488 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1217
timestamp 1435914306
transform 1 0 7488 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1218
timestamp 1435914306
transform 1 0 7488 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1219
timestamp 1435914306
transform 1 0 7488 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1220
timestamp 1435914306
transform 1 0 7488 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1221
timestamp 1435914306
transform 1 0 7488 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1222
timestamp 1435914306
transform 1 0 7488 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1223
timestamp 1435914306
transform 1 0 7488 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1224
timestamp 1435914306
transform 1 0 7488 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1225
timestamp 1435914306
transform 1 0 7488 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1226
timestamp 1435914306
transform 1 0 7488 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1227
timestamp 1435914306
transform 1 0 7488 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1228
timestamp 1435914306
transform 1 0 7488 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1229
timestamp 1435914306
transform 1 0 7488 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1230
timestamp 1435914306
transform 1 0 7488 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1231
timestamp 1435914306
transform 1 0 7488 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1232
timestamp 1435914306
transform 1 0 7488 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1233
timestamp 1435914306
transform 1 0 7488 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1234
timestamp 1435914306
transform 1 0 7488 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1235
timestamp 1435914306
transform 1 0 7488 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1236
timestamp 1435914306
transform 1 0 7488 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1237
timestamp 1435914306
transform 1 0 7488 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1238
timestamp 1435914306
transform 1 0 7488 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1239
timestamp 1435914306
transform 1 0 7488 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1240
timestamp 1435914306
transform 1 0 7488 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1241
timestamp 1435914306
transform 1 0 7488 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1242
timestamp 1435914306
transform 1 0 7488 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1243
timestamp 1435914306
transform 1 0 7488 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1244
timestamp 1435914306
transform 1 0 7488 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1245
timestamp 1435914306
transform 1 0 7488 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1246
timestamp 1435914306
transform 1 0 7488 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1247
timestamp 1435914306
transform 1 0 7488 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1248
timestamp 1435914306
transform 1 0 7488 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1249
timestamp 1435914306
transform 1 0 7488 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1250
timestamp 1435914306
transform 1 0 7488 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1251
timestamp 1435914306
transform 1 0 7488 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1252
timestamp 1435914306
transform 1 0 7488 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1253
timestamp 1435914306
transform 1 0 7488 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1254
timestamp 1435914306
transform 1 0 7488 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1255
timestamp 1435914306
transform 1 0 7488 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1256
timestamp 1435914306
transform 1 0 7488 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1257
timestamp 1435914306
transform 1 0 7488 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1258
timestamp 1435914306
transform 1 0 7488 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1259
timestamp 1435914306
transform 1 0 7488 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1260
timestamp 1435914306
transform 1 0 7488 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1261
timestamp 1435914306
transform 1 0 7488 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1262
timestamp 1435914306
transform 1 0 7488 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1263
timestamp 1435914306
transform 1 0 7488 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1264
timestamp 1435914306
transform 1 0 7488 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1265
timestamp 1435914306
transform 1 0 7488 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1266
timestamp 1435914306
transform 1 0 7488 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1267
timestamp 1435914306
transform 1 0 7488 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1268
timestamp 1435914306
transform 1 0 7488 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1269
timestamp 1435914306
transform 1 0 7488 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1270
timestamp 1435914306
transform 1 0 7488 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1271
timestamp 1435914306
transform 1 0 7488 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1272
timestamp 1435914306
transform 1 0 7488 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1273
timestamp 1435914306
transform 1 0 7488 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1274
timestamp 1435914306
transform 1 0 7488 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1275
timestamp 1435914306
transform 1 0 7488 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1276
timestamp 1435914306
transform 1 0 7488 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1277
timestamp 1435914306
transform 1 0 7488 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1278
timestamp 1435914306
transform 1 0 7488 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1279
timestamp 1435914306
transform 1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1280
timestamp 1435914306
transform -1 0 7488 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1281
timestamp 1435914306
transform -1 0 7488 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1282
timestamp 1435914306
transform -1 0 7488 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1283
timestamp 1435914306
transform -1 0 7488 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1284
timestamp 1435914306
transform -1 0 7488 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1285
timestamp 1435914306
transform -1 0 7488 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1286
timestamp 1435914306
transform -1 0 7488 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1287
timestamp 1435914306
transform -1 0 7488 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1288
timestamp 1435914306
transform -1 0 7488 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1289
timestamp 1435914306
transform -1 0 7488 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1290
timestamp 1435914306
transform -1 0 7488 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1291
timestamp 1435914306
transform -1 0 7488 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1292
timestamp 1435914306
transform -1 0 7488 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1293
timestamp 1435914306
transform -1 0 7488 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1294
timestamp 1435914306
transform -1 0 7488 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1295
timestamp 1435914306
transform -1 0 7488 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1296
timestamp 1435914306
transform -1 0 7488 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1297
timestamp 1435914306
transform -1 0 7488 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1298
timestamp 1435914306
transform -1 0 7488 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1299
timestamp 1435914306
transform -1 0 7488 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1300
timestamp 1435914306
transform -1 0 7488 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1301
timestamp 1435914306
transform -1 0 7488 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1302
timestamp 1435914306
transform -1 0 7488 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1303
timestamp 1435914306
transform -1 0 7488 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1304
timestamp 1435914306
transform -1 0 7488 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1305
timestamp 1435914306
transform -1 0 7488 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1306
timestamp 1435914306
transform -1 0 7488 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1307
timestamp 1435914306
transform -1 0 7488 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1308
timestamp 1435914306
transform -1 0 7488 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1309
timestamp 1435914306
transform -1 0 7488 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1310
timestamp 1435914306
transform -1 0 7488 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1311
timestamp 1435914306
transform -1 0 7488 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1312
timestamp 1435914306
transform -1 0 7488 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1313
timestamp 1435914306
transform -1 0 7488 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1314
timestamp 1435914306
transform -1 0 7488 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1315
timestamp 1435914306
transform -1 0 7488 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1316
timestamp 1435914306
transform -1 0 7488 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1317
timestamp 1435914306
transform -1 0 7488 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1318
timestamp 1435914306
transform -1 0 7488 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1319
timestamp 1435914306
transform -1 0 7488 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1320
timestamp 1435914306
transform -1 0 7488 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1321
timestamp 1435914306
transform -1 0 7488 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1322
timestamp 1435914306
transform -1 0 7488 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1323
timestamp 1435914306
transform -1 0 7488 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1324
timestamp 1435914306
transform -1 0 7488 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1325
timestamp 1435914306
transform -1 0 7488 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1326
timestamp 1435914306
transform -1 0 7488 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1327
timestamp 1435914306
transform -1 0 7488 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1328
timestamp 1435914306
transform -1 0 7488 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1329
timestamp 1435914306
transform -1 0 7488 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1330
timestamp 1435914306
transform -1 0 7488 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1331
timestamp 1435914306
transform -1 0 7488 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1332
timestamp 1435914306
transform -1 0 7488 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1333
timestamp 1435914306
transform -1 0 7488 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1334
timestamp 1435914306
transform -1 0 7488 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1335
timestamp 1435914306
transform -1 0 7488 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1336
timestamp 1435914306
transform -1 0 7488 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1337
timestamp 1435914306
transform -1 0 7488 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1338
timestamp 1435914306
transform -1 0 7488 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1339
timestamp 1435914306
transform -1 0 7488 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1340
timestamp 1435914306
transform -1 0 7488 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1341
timestamp 1435914306
transform -1 0 7488 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1342
timestamp 1435914306
transform -1 0 7488 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1343
timestamp 1435914306
transform -1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1344
timestamp 1435914306
transform 1 0 6240 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1345
timestamp 1435914306
transform 1 0 6240 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1346
timestamp 1435914306
transform 1 0 6240 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1347
timestamp 1435914306
transform 1 0 6240 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1348
timestamp 1435914306
transform 1 0 6240 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1349
timestamp 1435914306
transform 1 0 6240 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1350
timestamp 1435914306
transform 1 0 6240 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1351
timestamp 1435914306
transform 1 0 6240 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1352
timestamp 1435914306
transform 1 0 6240 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1353
timestamp 1435914306
transform 1 0 6240 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1354
timestamp 1435914306
transform 1 0 6240 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1355
timestamp 1435914306
transform 1 0 6240 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1356
timestamp 1435914306
transform 1 0 6240 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1357
timestamp 1435914306
transform 1 0 6240 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1358
timestamp 1435914306
transform 1 0 6240 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1359
timestamp 1435914306
transform 1 0 6240 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1360
timestamp 1435914306
transform 1 0 6240 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1361
timestamp 1435914306
transform 1 0 6240 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1362
timestamp 1435914306
transform 1 0 6240 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1363
timestamp 1435914306
transform 1 0 6240 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1364
timestamp 1435914306
transform 1 0 6240 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1365
timestamp 1435914306
transform 1 0 6240 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1366
timestamp 1435914306
transform 1 0 6240 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1367
timestamp 1435914306
transform 1 0 6240 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1368
timestamp 1435914306
transform 1 0 6240 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1369
timestamp 1435914306
transform 1 0 6240 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1370
timestamp 1435914306
transform 1 0 6240 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1371
timestamp 1435914306
transform 1 0 6240 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1372
timestamp 1435914306
transform 1 0 6240 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1373
timestamp 1435914306
transform 1 0 6240 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1374
timestamp 1435914306
transform 1 0 6240 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1375
timestamp 1435914306
transform 1 0 6240 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1376
timestamp 1435914306
transform 1 0 6240 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1377
timestamp 1435914306
transform 1 0 6240 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1378
timestamp 1435914306
transform 1 0 6240 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1379
timestamp 1435914306
transform 1 0 6240 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1380
timestamp 1435914306
transform 1 0 6240 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1381
timestamp 1435914306
transform 1 0 6240 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1382
timestamp 1435914306
transform 1 0 6240 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1383
timestamp 1435914306
transform 1 0 6240 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1384
timestamp 1435914306
transform 1 0 6240 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1385
timestamp 1435914306
transform 1 0 6240 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1386
timestamp 1435914306
transform 1 0 6240 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1387
timestamp 1435914306
transform 1 0 6240 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1388
timestamp 1435914306
transform 1 0 6240 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1389
timestamp 1435914306
transform 1 0 6240 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1390
timestamp 1435914306
transform 1 0 6240 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1391
timestamp 1435914306
transform 1 0 6240 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1392
timestamp 1435914306
transform 1 0 6240 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1393
timestamp 1435914306
transform 1 0 6240 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1394
timestamp 1435914306
transform 1 0 6240 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1395
timestamp 1435914306
transform 1 0 6240 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1396
timestamp 1435914306
transform 1 0 6240 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1397
timestamp 1435914306
transform 1 0 6240 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1398
timestamp 1435914306
transform 1 0 6240 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1399
timestamp 1435914306
transform 1 0 6240 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1400
timestamp 1435914306
transform 1 0 6240 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1401
timestamp 1435914306
transform 1 0 6240 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1402
timestamp 1435914306
transform 1 0 6240 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1403
timestamp 1435914306
transform 1 0 6240 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1404
timestamp 1435914306
transform 1 0 6240 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1405
timestamp 1435914306
transform 1 0 6240 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1406
timestamp 1435914306
transform 1 0 6240 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1407
timestamp 1435914306
transform 1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1408
timestamp 1435914306
transform -1 0 6240 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1409
timestamp 1435914306
transform -1 0 6240 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1410
timestamp 1435914306
transform -1 0 6240 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1411
timestamp 1435914306
transform -1 0 6240 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1412
timestamp 1435914306
transform -1 0 6240 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1413
timestamp 1435914306
transform -1 0 6240 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1414
timestamp 1435914306
transform -1 0 6240 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1415
timestamp 1435914306
transform -1 0 6240 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1416
timestamp 1435914306
transform -1 0 6240 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1417
timestamp 1435914306
transform -1 0 6240 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1418
timestamp 1435914306
transform -1 0 6240 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1419
timestamp 1435914306
transform -1 0 6240 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1420
timestamp 1435914306
transform -1 0 6240 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1421
timestamp 1435914306
transform -1 0 6240 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1422
timestamp 1435914306
transform -1 0 6240 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1423
timestamp 1435914306
transform -1 0 6240 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1424
timestamp 1435914306
transform -1 0 6240 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1425
timestamp 1435914306
transform -1 0 6240 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1426
timestamp 1435914306
transform -1 0 6240 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1427
timestamp 1435914306
transform -1 0 6240 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1428
timestamp 1435914306
transform -1 0 6240 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1429
timestamp 1435914306
transform -1 0 6240 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1430
timestamp 1435914306
transform -1 0 6240 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1431
timestamp 1435914306
transform -1 0 6240 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1432
timestamp 1435914306
transform -1 0 6240 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1433
timestamp 1435914306
transform -1 0 6240 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1434
timestamp 1435914306
transform -1 0 6240 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1435
timestamp 1435914306
transform -1 0 6240 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1436
timestamp 1435914306
transform -1 0 6240 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1437
timestamp 1435914306
transform -1 0 6240 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1438
timestamp 1435914306
transform -1 0 6240 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1439
timestamp 1435914306
transform -1 0 6240 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1440
timestamp 1435914306
transform -1 0 6240 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1441
timestamp 1435914306
transform -1 0 6240 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1442
timestamp 1435914306
transform -1 0 6240 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1443
timestamp 1435914306
transform -1 0 6240 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1444
timestamp 1435914306
transform -1 0 6240 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1445
timestamp 1435914306
transform -1 0 6240 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1446
timestamp 1435914306
transform -1 0 6240 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1447
timestamp 1435914306
transform -1 0 6240 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1448
timestamp 1435914306
transform -1 0 6240 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1449
timestamp 1435914306
transform -1 0 6240 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1450
timestamp 1435914306
transform -1 0 6240 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1451
timestamp 1435914306
transform -1 0 6240 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1452
timestamp 1435914306
transform -1 0 6240 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1453
timestamp 1435914306
transform -1 0 6240 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1454
timestamp 1435914306
transform -1 0 6240 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1455
timestamp 1435914306
transform -1 0 6240 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1456
timestamp 1435914306
transform -1 0 6240 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1457
timestamp 1435914306
transform -1 0 6240 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1458
timestamp 1435914306
transform -1 0 6240 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1459
timestamp 1435914306
transform -1 0 6240 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1460
timestamp 1435914306
transform -1 0 6240 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1461
timestamp 1435914306
transform -1 0 6240 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1462
timestamp 1435914306
transform -1 0 6240 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1463
timestamp 1435914306
transform -1 0 6240 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1464
timestamp 1435914306
transform -1 0 6240 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1465
timestamp 1435914306
transform -1 0 6240 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1466
timestamp 1435914306
transform -1 0 6240 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1467
timestamp 1435914306
transform -1 0 6240 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1468
timestamp 1435914306
transform -1 0 6240 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1469
timestamp 1435914306
transform -1 0 6240 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1470
timestamp 1435914306
transform -1 0 6240 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1471
timestamp 1435914306
transform -1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1472
timestamp 1435914306
transform 1 0 4992 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1473
timestamp 1435914306
transform 1 0 4992 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1474
timestamp 1435914306
transform 1 0 4992 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1475
timestamp 1435914306
transform 1 0 4992 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1476
timestamp 1435914306
transform 1 0 4992 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1477
timestamp 1435914306
transform 1 0 4992 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1478
timestamp 1435914306
transform 1 0 4992 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1479
timestamp 1435914306
transform 1 0 4992 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1480
timestamp 1435914306
transform 1 0 4992 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1481
timestamp 1435914306
transform 1 0 4992 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1482
timestamp 1435914306
transform 1 0 4992 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1483
timestamp 1435914306
transform 1 0 4992 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1484
timestamp 1435914306
transform 1 0 4992 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1485
timestamp 1435914306
transform 1 0 4992 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1486
timestamp 1435914306
transform 1 0 4992 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1487
timestamp 1435914306
transform 1 0 4992 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1488
timestamp 1435914306
transform 1 0 4992 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1489
timestamp 1435914306
transform 1 0 4992 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1490
timestamp 1435914306
transform 1 0 4992 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1491
timestamp 1435914306
transform 1 0 4992 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1492
timestamp 1435914306
transform 1 0 4992 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1493
timestamp 1435914306
transform 1 0 4992 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1494
timestamp 1435914306
transform 1 0 4992 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1495
timestamp 1435914306
transform 1 0 4992 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1496
timestamp 1435914306
transform 1 0 4992 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1497
timestamp 1435914306
transform 1 0 4992 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1498
timestamp 1435914306
transform 1 0 4992 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1499
timestamp 1435914306
transform 1 0 4992 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1500
timestamp 1435914306
transform 1 0 4992 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1501
timestamp 1435914306
transform 1 0 4992 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1502
timestamp 1435914306
transform 1 0 4992 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1503
timestamp 1435914306
transform 1 0 4992 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1504
timestamp 1435914306
transform 1 0 4992 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1505
timestamp 1435914306
transform 1 0 4992 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1506
timestamp 1435914306
transform 1 0 4992 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1507
timestamp 1435914306
transform 1 0 4992 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1508
timestamp 1435914306
transform 1 0 4992 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1509
timestamp 1435914306
transform 1 0 4992 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1510
timestamp 1435914306
transform 1 0 4992 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1511
timestamp 1435914306
transform 1 0 4992 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1512
timestamp 1435914306
transform 1 0 4992 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1513
timestamp 1435914306
transform 1 0 4992 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1514
timestamp 1435914306
transform 1 0 4992 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1515
timestamp 1435914306
transform 1 0 4992 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1516
timestamp 1435914306
transform 1 0 4992 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1517
timestamp 1435914306
transform 1 0 4992 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1518
timestamp 1435914306
transform 1 0 4992 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1519
timestamp 1435914306
transform 1 0 4992 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1520
timestamp 1435914306
transform 1 0 4992 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1521
timestamp 1435914306
transform 1 0 4992 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1522
timestamp 1435914306
transform 1 0 4992 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1523
timestamp 1435914306
transform 1 0 4992 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1524
timestamp 1435914306
transform 1 0 4992 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1525
timestamp 1435914306
transform 1 0 4992 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1526
timestamp 1435914306
transform 1 0 4992 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1527
timestamp 1435914306
transform 1 0 4992 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1528
timestamp 1435914306
transform 1 0 4992 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1529
timestamp 1435914306
transform 1 0 4992 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1530
timestamp 1435914306
transform 1 0 4992 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1531
timestamp 1435914306
transform 1 0 4992 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1532
timestamp 1435914306
transform 1 0 4992 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1533
timestamp 1435914306
transform 1 0 4992 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1534
timestamp 1435914306
transform 1 0 4992 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1535
timestamp 1435914306
transform 1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1536
timestamp 1435914306
transform -1 0 4992 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1537
timestamp 1435914306
transform -1 0 4992 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1538
timestamp 1435914306
transform -1 0 4992 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1539
timestamp 1435914306
transform -1 0 4992 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1540
timestamp 1435914306
transform -1 0 4992 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1541
timestamp 1435914306
transform -1 0 4992 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1542
timestamp 1435914306
transform -1 0 4992 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1543
timestamp 1435914306
transform -1 0 4992 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1544
timestamp 1435914306
transform -1 0 4992 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1545
timestamp 1435914306
transform -1 0 4992 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1546
timestamp 1435914306
transform -1 0 4992 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1547
timestamp 1435914306
transform -1 0 4992 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1548
timestamp 1435914306
transform -1 0 4992 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1549
timestamp 1435914306
transform -1 0 4992 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1550
timestamp 1435914306
transform -1 0 4992 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1551
timestamp 1435914306
transform -1 0 4992 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1552
timestamp 1435914306
transform -1 0 4992 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1553
timestamp 1435914306
transform -1 0 4992 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1554
timestamp 1435914306
transform -1 0 4992 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1555
timestamp 1435914306
transform -1 0 4992 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1556
timestamp 1435914306
transform -1 0 4992 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1557
timestamp 1435914306
transform -1 0 4992 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1558
timestamp 1435914306
transform -1 0 4992 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1559
timestamp 1435914306
transform -1 0 4992 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1560
timestamp 1435914306
transform -1 0 4992 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1561
timestamp 1435914306
transform -1 0 4992 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1562
timestamp 1435914306
transform -1 0 4992 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1563
timestamp 1435914306
transform -1 0 4992 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1564
timestamp 1435914306
transform -1 0 4992 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1565
timestamp 1435914306
transform -1 0 4992 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1566
timestamp 1435914306
transform -1 0 4992 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1567
timestamp 1435914306
transform -1 0 4992 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1568
timestamp 1435914306
transform -1 0 4992 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1569
timestamp 1435914306
transform -1 0 4992 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1570
timestamp 1435914306
transform -1 0 4992 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1571
timestamp 1435914306
transform -1 0 4992 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1572
timestamp 1435914306
transform -1 0 4992 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1573
timestamp 1435914306
transform -1 0 4992 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1574
timestamp 1435914306
transform -1 0 4992 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1575
timestamp 1435914306
transform -1 0 4992 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1576
timestamp 1435914306
transform -1 0 4992 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1577
timestamp 1435914306
transform -1 0 4992 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1578
timestamp 1435914306
transform -1 0 4992 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1579
timestamp 1435914306
transform -1 0 4992 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1580
timestamp 1435914306
transform -1 0 4992 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1581
timestamp 1435914306
transform -1 0 4992 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1582
timestamp 1435914306
transform -1 0 4992 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1583
timestamp 1435914306
transform -1 0 4992 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1584
timestamp 1435914306
transform -1 0 4992 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1585
timestamp 1435914306
transform -1 0 4992 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1586
timestamp 1435914306
transform -1 0 4992 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1587
timestamp 1435914306
transform -1 0 4992 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1588
timestamp 1435914306
transform -1 0 4992 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1589
timestamp 1435914306
transform -1 0 4992 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1590
timestamp 1435914306
transform -1 0 4992 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1591
timestamp 1435914306
transform -1 0 4992 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1592
timestamp 1435914306
transform -1 0 4992 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1593
timestamp 1435914306
transform -1 0 4992 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1594
timestamp 1435914306
transform -1 0 4992 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1595
timestamp 1435914306
transform -1 0 4992 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1596
timestamp 1435914306
transform -1 0 4992 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1597
timestamp 1435914306
transform -1 0 4992 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1598
timestamp 1435914306
transform -1 0 4992 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1599
timestamp 1435914306
transform -1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1600
timestamp 1435914306
transform 1 0 3744 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1601
timestamp 1435914306
transform 1 0 3744 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1602
timestamp 1435914306
transform 1 0 3744 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1603
timestamp 1435914306
transform 1 0 3744 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1604
timestamp 1435914306
transform 1 0 3744 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1605
timestamp 1435914306
transform 1 0 3744 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1606
timestamp 1435914306
transform 1 0 3744 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1607
timestamp 1435914306
transform 1 0 3744 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1608
timestamp 1435914306
transform 1 0 3744 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1609
timestamp 1435914306
transform 1 0 3744 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1610
timestamp 1435914306
transform 1 0 3744 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1611
timestamp 1435914306
transform 1 0 3744 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1612
timestamp 1435914306
transform 1 0 3744 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1613
timestamp 1435914306
transform 1 0 3744 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1614
timestamp 1435914306
transform 1 0 3744 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1615
timestamp 1435914306
transform 1 0 3744 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1616
timestamp 1435914306
transform 1 0 3744 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1617
timestamp 1435914306
transform 1 0 3744 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1618
timestamp 1435914306
transform 1 0 3744 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1619
timestamp 1435914306
transform 1 0 3744 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1620
timestamp 1435914306
transform 1 0 3744 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1621
timestamp 1435914306
transform 1 0 3744 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1622
timestamp 1435914306
transform 1 0 3744 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1623
timestamp 1435914306
transform 1 0 3744 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1624
timestamp 1435914306
transform 1 0 3744 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1625
timestamp 1435914306
transform 1 0 3744 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1626
timestamp 1435914306
transform 1 0 3744 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1627
timestamp 1435914306
transform 1 0 3744 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1628
timestamp 1435914306
transform 1 0 3744 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1629
timestamp 1435914306
transform 1 0 3744 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1630
timestamp 1435914306
transform 1 0 3744 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1631
timestamp 1435914306
transform 1 0 3744 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1632
timestamp 1435914306
transform 1 0 3744 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1633
timestamp 1435914306
transform 1 0 3744 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1634
timestamp 1435914306
transform 1 0 3744 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1635
timestamp 1435914306
transform 1 0 3744 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1636
timestamp 1435914306
transform 1 0 3744 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1637
timestamp 1435914306
transform 1 0 3744 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1638
timestamp 1435914306
transform 1 0 3744 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1639
timestamp 1435914306
transform 1 0 3744 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1640
timestamp 1435914306
transform 1 0 3744 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1641
timestamp 1435914306
transform 1 0 3744 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1642
timestamp 1435914306
transform 1 0 3744 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1643
timestamp 1435914306
transform 1 0 3744 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1644
timestamp 1435914306
transform 1 0 3744 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1645
timestamp 1435914306
transform 1 0 3744 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1646
timestamp 1435914306
transform 1 0 3744 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1647
timestamp 1435914306
transform 1 0 3744 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1648
timestamp 1435914306
transform 1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1649
timestamp 1435914306
transform 1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1650
timestamp 1435914306
transform 1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1651
timestamp 1435914306
transform 1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1652
timestamp 1435914306
transform 1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1653
timestamp 1435914306
transform 1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1654
timestamp 1435914306
transform 1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1655
timestamp 1435914306
transform 1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1656
timestamp 1435914306
transform 1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1657
timestamp 1435914306
transform 1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1658
timestamp 1435914306
transform 1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1659
timestamp 1435914306
transform 1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1660
timestamp 1435914306
transform 1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1661
timestamp 1435914306
transform 1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1662
timestamp 1435914306
transform 1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1663
timestamp 1435914306
transform 1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1664
timestamp 1435914306
transform -1 0 3744 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1665
timestamp 1435914306
transform -1 0 3744 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1666
timestamp 1435914306
transform -1 0 3744 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1667
timestamp 1435914306
transform -1 0 3744 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1668
timestamp 1435914306
transform -1 0 3744 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1669
timestamp 1435914306
transform -1 0 3744 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1670
timestamp 1435914306
transform -1 0 3744 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1671
timestamp 1435914306
transform -1 0 3744 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1672
timestamp 1435914306
transform -1 0 3744 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1673
timestamp 1435914306
transform -1 0 3744 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1674
timestamp 1435914306
transform -1 0 3744 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1675
timestamp 1435914306
transform -1 0 3744 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1676
timestamp 1435914306
transform -1 0 3744 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1677
timestamp 1435914306
transform -1 0 3744 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1678
timestamp 1435914306
transform -1 0 3744 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1679
timestamp 1435914306
transform -1 0 3744 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1680
timestamp 1435914306
transform -1 0 3744 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1681
timestamp 1435914306
transform -1 0 3744 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1682
timestamp 1435914306
transform -1 0 3744 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1683
timestamp 1435914306
transform -1 0 3744 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1684
timestamp 1435914306
transform -1 0 3744 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1685
timestamp 1435914306
transform -1 0 3744 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1686
timestamp 1435914306
transform -1 0 3744 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1687
timestamp 1435914306
transform -1 0 3744 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1688
timestamp 1435914306
transform -1 0 3744 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1689
timestamp 1435914306
transform -1 0 3744 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1690
timestamp 1435914306
transform -1 0 3744 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1691
timestamp 1435914306
transform -1 0 3744 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1692
timestamp 1435914306
transform -1 0 3744 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1693
timestamp 1435914306
transform -1 0 3744 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1694
timestamp 1435914306
transform -1 0 3744 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1695
timestamp 1435914306
transform -1 0 3744 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1696
timestamp 1435914306
transform -1 0 3744 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1697
timestamp 1435914306
transform -1 0 3744 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1698
timestamp 1435914306
transform -1 0 3744 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1699
timestamp 1435914306
transform -1 0 3744 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1700
timestamp 1435914306
transform -1 0 3744 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1701
timestamp 1435914306
transform -1 0 3744 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1702
timestamp 1435914306
transform -1 0 3744 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1703
timestamp 1435914306
transform -1 0 3744 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1704
timestamp 1435914306
transform -1 0 3744 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1705
timestamp 1435914306
transform -1 0 3744 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1706
timestamp 1435914306
transform -1 0 3744 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1707
timestamp 1435914306
transform -1 0 3744 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1708
timestamp 1435914306
transform -1 0 3744 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1709
timestamp 1435914306
transform -1 0 3744 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1710
timestamp 1435914306
transform -1 0 3744 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1711
timestamp 1435914306
transform -1 0 3744 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1712
timestamp 1435914306
transform -1 0 3744 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1713
timestamp 1435914306
transform -1 0 3744 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1714
timestamp 1435914306
transform -1 0 3744 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1715
timestamp 1435914306
transform -1 0 3744 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1716
timestamp 1435914306
transform -1 0 3744 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1717
timestamp 1435914306
transform -1 0 3744 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1718
timestamp 1435914306
transform -1 0 3744 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1719
timestamp 1435914306
transform -1 0 3744 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1720
timestamp 1435914306
transform -1 0 3744 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1721
timestamp 1435914306
transform -1 0 3744 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1722
timestamp 1435914306
transform -1 0 3744 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1723
timestamp 1435914306
transform -1 0 3744 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1724
timestamp 1435914306
transform -1 0 3744 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1725
timestamp 1435914306
transform -1 0 3744 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1726
timestamp 1435914306
transform -1 0 3744 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1727
timestamp 1435914306
transform -1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1728
timestamp 1435914306
transform 1 0 2496 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1729
timestamp 1435914306
transform 1 0 2496 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1730
timestamp 1435914306
transform 1 0 2496 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1731
timestamp 1435914306
transform 1 0 2496 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1732
timestamp 1435914306
transform 1 0 2496 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1733
timestamp 1435914306
transform 1 0 2496 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1734
timestamp 1435914306
transform 1 0 2496 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1735
timestamp 1435914306
transform 1 0 2496 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1736
timestamp 1435914306
transform 1 0 2496 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1737
timestamp 1435914306
transform 1 0 2496 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1738
timestamp 1435914306
transform 1 0 2496 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1739
timestamp 1435914306
transform 1 0 2496 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1740
timestamp 1435914306
transform 1 0 2496 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1741
timestamp 1435914306
transform 1 0 2496 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1742
timestamp 1435914306
transform 1 0 2496 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1743
timestamp 1435914306
transform 1 0 2496 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1744
timestamp 1435914306
transform 1 0 2496 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1745
timestamp 1435914306
transform 1 0 2496 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1746
timestamp 1435914306
transform 1 0 2496 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1747
timestamp 1435914306
transform 1 0 2496 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1748
timestamp 1435914306
transform 1 0 2496 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1749
timestamp 1435914306
transform 1 0 2496 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1750
timestamp 1435914306
transform 1 0 2496 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1751
timestamp 1435914306
transform 1 0 2496 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1752
timestamp 1435914306
transform 1 0 2496 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1753
timestamp 1435914306
transform 1 0 2496 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1754
timestamp 1435914306
transform 1 0 2496 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1755
timestamp 1435914306
transform 1 0 2496 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1756
timestamp 1435914306
transform 1 0 2496 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1757
timestamp 1435914306
transform 1 0 2496 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1758
timestamp 1435914306
transform 1 0 2496 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1759
timestamp 1435914306
transform 1 0 2496 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1760
timestamp 1435914306
transform 1 0 2496 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1761
timestamp 1435914306
transform 1 0 2496 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1762
timestamp 1435914306
transform 1 0 2496 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1763
timestamp 1435914306
transform 1 0 2496 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1764
timestamp 1435914306
transform 1 0 2496 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1765
timestamp 1435914306
transform 1 0 2496 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1766
timestamp 1435914306
transform 1 0 2496 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1767
timestamp 1435914306
transform 1 0 2496 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1768
timestamp 1435914306
transform 1 0 2496 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1769
timestamp 1435914306
transform 1 0 2496 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1770
timestamp 1435914306
transform 1 0 2496 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1771
timestamp 1435914306
transform 1 0 2496 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1772
timestamp 1435914306
transform 1 0 2496 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1773
timestamp 1435914306
transform 1 0 2496 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1774
timestamp 1435914306
transform 1 0 2496 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1775
timestamp 1435914306
transform 1 0 2496 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1776
timestamp 1435914306
transform 1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1777
timestamp 1435914306
transform 1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1778
timestamp 1435914306
transform 1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1779
timestamp 1435914306
transform 1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1780
timestamp 1435914306
transform 1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1781
timestamp 1435914306
transform 1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1782
timestamp 1435914306
transform 1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1783
timestamp 1435914306
transform 1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1784
timestamp 1435914306
transform 1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1785
timestamp 1435914306
transform 1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1786
timestamp 1435914306
transform 1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1787
timestamp 1435914306
transform 1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1788
timestamp 1435914306
transform 1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1789
timestamp 1435914306
transform 1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1790
timestamp 1435914306
transform 1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1791
timestamp 1435914306
transform 1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1792
timestamp 1435914306
transform -1 0 2496 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1793
timestamp 1435914306
transform -1 0 2496 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1794
timestamp 1435914306
transform -1 0 2496 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1795
timestamp 1435914306
transform -1 0 2496 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1796
timestamp 1435914306
transform -1 0 2496 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1797
timestamp 1435914306
transform -1 0 2496 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1798
timestamp 1435914306
transform -1 0 2496 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1799
timestamp 1435914306
transform -1 0 2496 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1800
timestamp 1435914306
transform -1 0 2496 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1801
timestamp 1435914306
transform -1 0 2496 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1802
timestamp 1435914306
transform -1 0 2496 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1803
timestamp 1435914306
transform -1 0 2496 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1804
timestamp 1435914306
transform -1 0 2496 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1805
timestamp 1435914306
transform -1 0 2496 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1806
timestamp 1435914306
transform -1 0 2496 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1807
timestamp 1435914306
transform -1 0 2496 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1808
timestamp 1435914306
transform -1 0 2496 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1809
timestamp 1435914306
transform -1 0 2496 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1810
timestamp 1435914306
transform -1 0 2496 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1811
timestamp 1435914306
transform -1 0 2496 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1812
timestamp 1435914306
transform -1 0 2496 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1813
timestamp 1435914306
transform -1 0 2496 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1814
timestamp 1435914306
transform -1 0 2496 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1815
timestamp 1435914306
transform -1 0 2496 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1816
timestamp 1435914306
transform -1 0 2496 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1817
timestamp 1435914306
transform -1 0 2496 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1818
timestamp 1435914306
transform -1 0 2496 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1819
timestamp 1435914306
transform -1 0 2496 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1820
timestamp 1435914306
transform -1 0 2496 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1821
timestamp 1435914306
transform -1 0 2496 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1822
timestamp 1435914306
transform -1 0 2496 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1823
timestamp 1435914306
transform -1 0 2496 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1824
timestamp 1435914306
transform -1 0 2496 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1825
timestamp 1435914306
transform -1 0 2496 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1826
timestamp 1435914306
transform -1 0 2496 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1827
timestamp 1435914306
transform -1 0 2496 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1828
timestamp 1435914306
transform -1 0 2496 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1829
timestamp 1435914306
transform -1 0 2496 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1830
timestamp 1435914306
transform -1 0 2496 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1831
timestamp 1435914306
transform -1 0 2496 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1832
timestamp 1435914306
transform -1 0 2496 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1833
timestamp 1435914306
transform -1 0 2496 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1834
timestamp 1435914306
transform -1 0 2496 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1835
timestamp 1435914306
transform -1 0 2496 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1836
timestamp 1435914306
transform -1 0 2496 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1837
timestamp 1435914306
transform -1 0 2496 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1838
timestamp 1435914306
transform -1 0 2496 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1839
timestamp 1435914306
transform -1 0 2496 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1840
timestamp 1435914306
transform -1 0 2496 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1841
timestamp 1435914306
transform -1 0 2496 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1842
timestamp 1435914306
transform -1 0 2496 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1843
timestamp 1435914306
transform -1 0 2496 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1844
timestamp 1435914306
transform -1 0 2496 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1845
timestamp 1435914306
transform -1 0 2496 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1846
timestamp 1435914306
transform -1 0 2496 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1847
timestamp 1435914306
transform -1 0 2496 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1848
timestamp 1435914306
transform -1 0 2496 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1849
timestamp 1435914306
transform -1 0 2496 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1850
timestamp 1435914306
transform -1 0 2496 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1851
timestamp 1435914306
transform -1 0 2496 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1852
timestamp 1435914306
transform -1 0 2496 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1853
timestamp 1435914306
transform -1 0 2496 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1854
timestamp 1435914306
transform -1 0 2496 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1855
timestamp 1435914306
transform -1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1856
timestamp 1435914306
transform 1 0 1248 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1857
timestamp 1435914306
transform 1 0 1248 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1858
timestamp 1435914306
transform 1 0 1248 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1859
timestamp 1435914306
transform 1 0 1248 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1860
timestamp 1435914306
transform 1 0 1248 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1861
timestamp 1435914306
transform 1 0 1248 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1862
timestamp 1435914306
transform 1 0 1248 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1863
timestamp 1435914306
transform 1 0 1248 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1864
timestamp 1435914306
transform 1 0 1248 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1865
timestamp 1435914306
transform 1 0 1248 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1866
timestamp 1435914306
transform 1 0 1248 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1867
timestamp 1435914306
transform 1 0 1248 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1868
timestamp 1435914306
transform 1 0 1248 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1869
timestamp 1435914306
transform 1 0 1248 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1870
timestamp 1435914306
transform 1 0 1248 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1871
timestamp 1435914306
transform 1 0 1248 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1872
timestamp 1435914306
transform 1 0 1248 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1873
timestamp 1435914306
transform 1 0 1248 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1874
timestamp 1435914306
transform 1 0 1248 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1875
timestamp 1435914306
transform 1 0 1248 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1876
timestamp 1435914306
transform 1 0 1248 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1877
timestamp 1435914306
transform 1 0 1248 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1878
timestamp 1435914306
transform 1 0 1248 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1879
timestamp 1435914306
transform 1 0 1248 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1880
timestamp 1435914306
transform 1 0 1248 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1881
timestamp 1435914306
transform 1 0 1248 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1882
timestamp 1435914306
transform 1 0 1248 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1883
timestamp 1435914306
transform 1 0 1248 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1884
timestamp 1435914306
transform 1 0 1248 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1885
timestamp 1435914306
transform 1 0 1248 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1886
timestamp 1435914306
transform 1 0 1248 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1887
timestamp 1435914306
transform 1 0 1248 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1888
timestamp 1435914306
transform 1 0 1248 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1889
timestamp 1435914306
transform 1 0 1248 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1890
timestamp 1435914306
transform 1 0 1248 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1891
timestamp 1435914306
transform 1 0 1248 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1892
timestamp 1435914306
transform 1 0 1248 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1893
timestamp 1435914306
transform 1 0 1248 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1894
timestamp 1435914306
transform 1 0 1248 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1895
timestamp 1435914306
transform 1 0 1248 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1896
timestamp 1435914306
transform 1 0 1248 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1897
timestamp 1435914306
transform 1 0 1248 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1898
timestamp 1435914306
transform 1 0 1248 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1899
timestamp 1435914306
transform 1 0 1248 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1900
timestamp 1435914306
transform 1 0 1248 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1901
timestamp 1435914306
transform 1 0 1248 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1902
timestamp 1435914306
transform 1 0 1248 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1903
timestamp 1435914306
transform 1 0 1248 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1904
timestamp 1435914306
transform 1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1905
timestamp 1435914306
transform 1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1906
timestamp 1435914306
transform 1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1907
timestamp 1435914306
transform 1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1908
timestamp 1435914306
transform 1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1909
timestamp 1435914306
transform 1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1910
timestamp 1435914306
transform 1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1911
timestamp 1435914306
transform 1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1912
timestamp 1435914306
transform 1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1913
timestamp 1435914306
transform 1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1914
timestamp 1435914306
transform 1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1915
timestamp 1435914306
transform 1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1916
timestamp 1435914306
transform 1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1917
timestamp 1435914306
transform 1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1918
timestamp 1435914306
transform 1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1919
timestamp 1435914306
transform 1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1920
timestamp 1435914306
transform -1 0 1248 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1921
timestamp 1435914306
transform -1 0 1248 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1922
timestamp 1435914306
transform -1 0 1248 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1923
timestamp 1435914306
transform -1 0 1248 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1924
timestamp 1435914306
transform -1 0 1248 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1925
timestamp 1435914306
transform -1 0 1248 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1926
timestamp 1435914306
transform -1 0 1248 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1927
timestamp 1435914306
transform -1 0 1248 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1928
timestamp 1435914306
transform -1 0 1248 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1929
timestamp 1435914306
transform -1 0 1248 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1930
timestamp 1435914306
transform -1 0 1248 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1931
timestamp 1435914306
transform -1 0 1248 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1932
timestamp 1435914306
transform -1 0 1248 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1933
timestamp 1435914306
transform -1 0 1248 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1934
timestamp 1435914306
transform -1 0 1248 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1935
timestamp 1435914306
transform -1 0 1248 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1936
timestamp 1435914306
transform -1 0 1248 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1937
timestamp 1435914306
transform -1 0 1248 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1938
timestamp 1435914306
transform -1 0 1248 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1939
timestamp 1435914306
transform -1 0 1248 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1940
timestamp 1435914306
transform -1 0 1248 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1941
timestamp 1435914306
transform -1 0 1248 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1942
timestamp 1435914306
transform -1 0 1248 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1943
timestamp 1435914306
transform -1 0 1248 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1944
timestamp 1435914306
transform -1 0 1248 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1945
timestamp 1435914306
transform -1 0 1248 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1946
timestamp 1435914306
transform -1 0 1248 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1947
timestamp 1435914306
transform -1 0 1248 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1948
timestamp 1435914306
transform -1 0 1248 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1949
timestamp 1435914306
transform -1 0 1248 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1950
timestamp 1435914306
transform -1 0 1248 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1951
timestamp 1435914306
transform -1 0 1248 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1952
timestamp 1435914306
transform -1 0 1248 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1953
timestamp 1435914306
transform -1 0 1248 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1954
timestamp 1435914306
transform -1 0 1248 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1955
timestamp 1435914306
transform -1 0 1248 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1956
timestamp 1435914306
transform -1 0 1248 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1957
timestamp 1435914306
transform -1 0 1248 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1958
timestamp 1435914306
transform -1 0 1248 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1959
timestamp 1435914306
transform -1 0 1248 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1960
timestamp 1435914306
transform -1 0 1248 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1961
timestamp 1435914306
transform -1 0 1248 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1962
timestamp 1435914306
transform -1 0 1248 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1963
timestamp 1435914306
transform -1 0 1248 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1964
timestamp 1435914306
transform -1 0 1248 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1965
timestamp 1435914306
transform -1 0 1248 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1966
timestamp 1435914306
transform -1 0 1248 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1967
timestamp 1435914306
transform -1 0 1248 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1968
timestamp 1435914306
transform -1 0 1248 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1969
timestamp 1435914306
transform -1 0 1248 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1970
timestamp 1435914306
transform -1 0 1248 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1971
timestamp 1435914306
transform -1 0 1248 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1972
timestamp 1435914306
transform -1 0 1248 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1973
timestamp 1435914306
transform -1 0 1248 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1974
timestamp 1435914306
transform -1 0 1248 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1975
timestamp 1435914306
transform -1 0 1248 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1976
timestamp 1435914306
transform -1 0 1248 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1977
timestamp 1435914306
transform -1 0 1248 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1978
timestamp 1435914306
transform -1 0 1248 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1979
timestamp 1435914306
transform -1 0 1248 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1980
timestamp 1435914306
transform -1 0 1248 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1981
timestamp 1435914306
transform -1 0 1248 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1982
timestamp 1435914306
transform -1 0 1248 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1983
timestamp 1435914306
transform -1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1984
timestamp 1435914306
transform 1 0 0 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1985
timestamp 1435914306
transform 1 0 0 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1986
timestamp 1435914306
transform 1 0 0 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1987
timestamp 1435914306
transform 1 0 0 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1988
timestamp 1435914306
transform 1 0 0 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1989
timestamp 1435914306
transform 1 0 0 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1990
timestamp 1435914306
transform 1 0 0 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1991
timestamp 1435914306
transform 1 0 0 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1992
timestamp 1435914306
transform 1 0 0 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1993
timestamp 1435914306
transform 1 0 0 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1994
timestamp 1435914306
transform 1 0 0 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1995
timestamp 1435914306
transform 1 0 0 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1996
timestamp 1435914306
transform 1 0 0 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1997
timestamp 1435914306
transform 1 0 0 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1998
timestamp 1435914306
transform 1 0 0 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_1999
timestamp 1435914306
transform 1 0 0 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2000
timestamp 1435914306
transform 1 0 0 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2001
timestamp 1435914306
transform 1 0 0 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2002
timestamp 1435914306
transform 1 0 0 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2003
timestamp 1435914306
transform 1 0 0 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2004
timestamp 1435914306
transform 1 0 0 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2005
timestamp 1435914306
transform 1 0 0 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2006
timestamp 1435914306
transform 1 0 0 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2007
timestamp 1435914306
transform 1 0 0 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2008
timestamp 1435914306
transform 1 0 0 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2009
timestamp 1435914306
transform 1 0 0 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2010
timestamp 1435914306
transform 1 0 0 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2011
timestamp 1435914306
transform 1 0 0 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2012
timestamp 1435914306
transform 1 0 0 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2013
timestamp 1435914306
transform 1 0 0 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2014
timestamp 1435914306
transform 1 0 0 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2015
timestamp 1435914306
transform 1 0 0 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2016
timestamp 1435914306
transform 1 0 0 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2017
timestamp 1435914306
transform 1 0 0 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2018
timestamp 1435914306
transform 1 0 0 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2019
timestamp 1435914306
transform 1 0 0 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2020
timestamp 1435914306
transform 1 0 0 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2021
timestamp 1435914306
transform 1 0 0 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2022
timestamp 1435914306
transform 1 0 0 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2023
timestamp 1435914306
transform 1 0 0 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2024
timestamp 1435914306
transform 1 0 0 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2025
timestamp 1435914306
transform 1 0 0 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2026
timestamp 1435914306
transform 1 0 0 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2027
timestamp 1435914306
transform 1 0 0 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2028
timestamp 1435914306
transform 1 0 0 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2029
timestamp 1435914306
transform 1 0 0 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2030
timestamp 1435914306
transform 1 0 0 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2031
timestamp 1435914306
transform 1 0 0 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2032
timestamp 1435914306
transform 1 0 0 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2033
timestamp 1435914306
transform 1 0 0 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2034
timestamp 1435914306
transform 1 0 0 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2035
timestamp 1435914306
transform 1 0 0 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2036
timestamp 1435914306
transform 1 0 0 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2037
timestamp 1435914306
transform 1 0 0 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2038
timestamp 1435914306
transform 1 0 0 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2039
timestamp 1435914306
transform 1 0 0 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2040
timestamp 1435914306
transform 1 0 0 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2041
timestamp 1435914306
transform 1 0 0 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2042
timestamp 1435914306
transform 1 0 0 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2043
timestamp 1435914306
transform 1 0 0 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2044
timestamp 1435914306
transform 1 0 0 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2045
timestamp 1435914306
transform 1 0 0 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2046
timestamp 1435914306
transform 1 0 0 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell  sky130_fd_bd_sram__openram_dp_cell_2047
timestamp 1435914306
transform 1 0 0 0 1 0
box -42 -105 650 421
<< labels >>
rlabel metal1 s 78 0 114 25280 4 bl_0_0
port 3 nsew
rlabel metal1 s 150 0 186 25280 4 br_0_0
port 5 nsew
rlabel metal1 s 294 0 330 25280 4 bl_1_0
port 7 nsew
rlabel metal1 s 366 0 402 25280 4 br_1_0
port 9 nsew
rlabel metal1 s 1134 0 1170 25280 4 bl_0_1
port 11 nsew
rlabel metal1 s 1062 0 1098 25280 4 br_0_1
port 13 nsew
rlabel metal1 s 918 0 954 25280 4 bl_1_1
port 15 nsew
rlabel metal1 s 846 0 882 25280 4 br_1_1
port 17 nsew
rlabel metal1 s 1326 0 1362 25280 4 bl_0_2
port 19 nsew
rlabel metal1 s 1398 0 1434 25280 4 br_0_2
port 21 nsew
rlabel metal1 s 1542 0 1578 25280 4 bl_1_2
port 23 nsew
rlabel metal1 s 1614 0 1650 25280 4 br_1_2
port 25 nsew
rlabel metal1 s 2382 0 2418 25280 4 bl_0_3
port 27 nsew
rlabel metal1 s 2310 0 2346 25280 4 br_0_3
port 29 nsew
rlabel metal1 s 2166 0 2202 25280 4 bl_1_3
port 31 nsew
rlabel metal1 s 2094 0 2130 25280 4 br_1_3
port 33 nsew
rlabel metal1 s 2574 0 2610 25280 4 bl_0_4
port 35 nsew
rlabel metal1 s 2646 0 2682 25280 4 br_0_4
port 37 nsew
rlabel metal1 s 2790 0 2826 25280 4 bl_1_4
port 39 nsew
rlabel metal1 s 2862 0 2898 25280 4 br_1_4
port 41 nsew
rlabel metal1 s 3630 0 3666 25280 4 bl_0_5
port 43 nsew
rlabel metal1 s 3558 0 3594 25280 4 br_0_5
port 45 nsew
rlabel metal1 s 3414 0 3450 25280 4 bl_1_5
port 47 nsew
rlabel metal1 s 3342 0 3378 25280 4 br_1_5
port 49 nsew
rlabel metal1 s 3822 0 3858 25280 4 bl_0_6
port 51 nsew
rlabel metal1 s 3894 0 3930 25280 4 br_0_6
port 53 nsew
rlabel metal1 s 4038 0 4074 25280 4 bl_1_6
port 55 nsew
rlabel metal1 s 4110 0 4146 25280 4 br_1_6
port 57 nsew
rlabel metal1 s 4878 0 4914 25280 4 bl_0_7
port 59 nsew
rlabel metal1 s 4806 0 4842 25280 4 br_0_7
port 61 nsew
rlabel metal1 s 4662 0 4698 25280 4 bl_1_7
port 63 nsew
rlabel metal1 s 4590 0 4626 25280 4 br_1_7
port 65 nsew
rlabel metal1 s 5070 0 5106 25280 4 bl_0_8
port 67 nsew
rlabel metal1 s 5142 0 5178 25280 4 br_0_8
port 69 nsew
rlabel metal1 s 5286 0 5322 25280 4 bl_1_8
port 71 nsew
rlabel metal1 s 5358 0 5394 25280 4 br_1_8
port 73 nsew
rlabel metal1 s 6126 0 6162 25280 4 bl_0_9
port 75 nsew
rlabel metal1 s 6054 0 6090 25280 4 br_0_9
port 77 nsew
rlabel metal1 s 5910 0 5946 25280 4 bl_1_9
port 79 nsew
rlabel metal1 s 5838 0 5874 25280 4 br_1_9
port 81 nsew
rlabel metal1 s 6318 0 6354 25280 4 bl_0_10
port 83 nsew
rlabel metal1 s 6390 0 6426 25280 4 br_0_10
port 85 nsew
rlabel metal1 s 6534 0 6570 25280 4 bl_1_10
port 87 nsew
rlabel metal1 s 6606 0 6642 25280 4 br_1_10
port 89 nsew
rlabel metal1 s 7374 0 7410 25280 4 bl_0_11
port 91 nsew
rlabel metal1 s 7302 0 7338 25280 4 br_0_11
port 93 nsew
rlabel metal1 s 7158 0 7194 25280 4 bl_1_11
port 95 nsew
rlabel metal1 s 7086 0 7122 25280 4 br_1_11
port 97 nsew
rlabel metal1 s 7566 0 7602 25280 4 bl_0_12
port 99 nsew
rlabel metal1 s 7638 0 7674 25280 4 br_0_12
port 101 nsew
rlabel metal1 s 7782 0 7818 25280 4 bl_1_12
port 103 nsew
rlabel metal1 s 7854 0 7890 25280 4 br_1_12
port 105 nsew
rlabel metal1 s 8622 0 8658 25280 4 bl_0_13
port 107 nsew
rlabel metal1 s 8550 0 8586 25280 4 br_0_13
port 109 nsew
rlabel metal1 s 8406 0 8442 25280 4 bl_1_13
port 111 nsew
rlabel metal1 s 8334 0 8370 25280 4 br_1_13
port 113 nsew
rlabel metal1 s 8814 0 8850 25280 4 bl_0_14
port 115 nsew
rlabel metal1 s 8886 0 8922 25280 4 br_0_14
port 117 nsew
rlabel metal1 s 9030 0 9066 25280 4 bl_1_14
port 119 nsew
rlabel metal1 s 9102 0 9138 25280 4 br_1_14
port 121 nsew
rlabel metal1 s 9870 0 9906 25280 4 bl_0_15
port 123 nsew
rlabel metal1 s 9798 0 9834 25280 4 br_0_15
port 125 nsew
rlabel metal1 s 9654 0 9690 25280 4 bl_1_15
port 127 nsew
rlabel metal1 s 9582 0 9618 25280 4 br_1_15
port 129 nsew
rlabel metal1 s 10062 0 10098 25280 4 bl_0_16
port 131 nsew
rlabel metal1 s 10134 0 10170 25280 4 br_0_16
port 133 nsew
rlabel metal1 s 10278 0 10314 25280 4 bl_1_16
port 135 nsew
rlabel metal1 s 10350 0 10386 25280 4 br_1_16
port 137 nsew
rlabel metal1 s 11118 0 11154 25280 4 bl_0_17
port 139 nsew
rlabel metal1 s 11046 0 11082 25280 4 br_0_17
port 141 nsew
rlabel metal1 s 10902 0 10938 25280 4 bl_1_17
port 143 nsew
rlabel metal1 s 10830 0 10866 25280 4 br_1_17
port 145 nsew
rlabel metal1 s 11310 0 11346 25280 4 bl_0_18
port 147 nsew
rlabel metal1 s 11382 0 11418 25280 4 br_0_18
port 149 nsew
rlabel metal1 s 11526 0 11562 25280 4 bl_1_18
port 151 nsew
rlabel metal1 s 11598 0 11634 25280 4 br_1_18
port 153 nsew
rlabel metal1 s 12366 0 12402 25280 4 bl_0_19
port 155 nsew
rlabel metal1 s 12294 0 12330 25280 4 br_0_19
port 157 nsew
rlabel metal1 s 12150 0 12186 25280 4 bl_1_19
port 159 nsew
rlabel metal1 s 12078 0 12114 25280 4 br_1_19
port 161 nsew
rlabel metal1 s 12558 0 12594 25280 4 bl_0_20
port 163 nsew
rlabel metal1 s 12630 0 12666 25280 4 br_0_20
port 165 nsew
rlabel metal1 s 12774 0 12810 25280 4 bl_1_20
port 167 nsew
rlabel metal1 s 12846 0 12882 25280 4 br_1_20
port 169 nsew
rlabel metal1 s 13614 0 13650 25280 4 bl_0_21
port 171 nsew
rlabel metal1 s 13542 0 13578 25280 4 br_0_21
port 173 nsew
rlabel metal1 s 13398 0 13434 25280 4 bl_1_21
port 175 nsew
rlabel metal1 s 13326 0 13362 25280 4 br_1_21
port 177 nsew
rlabel metal1 s 13806 0 13842 25280 4 bl_0_22
port 179 nsew
rlabel metal1 s 13878 0 13914 25280 4 br_0_22
port 181 nsew
rlabel metal1 s 14022 0 14058 25280 4 bl_1_22
port 183 nsew
rlabel metal1 s 14094 0 14130 25280 4 br_1_22
port 185 nsew
rlabel metal1 s 14862 0 14898 25280 4 bl_0_23
port 187 nsew
rlabel metal1 s 14790 0 14826 25280 4 br_0_23
port 189 nsew
rlabel metal1 s 14646 0 14682 25280 4 bl_1_23
port 191 nsew
rlabel metal1 s 14574 0 14610 25280 4 br_1_23
port 193 nsew
rlabel metal1 s 15054 0 15090 25280 4 bl_0_24
port 195 nsew
rlabel metal1 s 15126 0 15162 25280 4 br_0_24
port 197 nsew
rlabel metal1 s 15270 0 15306 25280 4 bl_1_24
port 199 nsew
rlabel metal1 s 15342 0 15378 25280 4 br_1_24
port 201 nsew
rlabel metal1 s 16110 0 16146 25280 4 bl_0_25
port 203 nsew
rlabel metal1 s 16038 0 16074 25280 4 br_0_25
port 205 nsew
rlabel metal1 s 15894 0 15930 25280 4 bl_1_25
port 207 nsew
rlabel metal1 s 15822 0 15858 25280 4 br_1_25
port 209 nsew
rlabel metal1 s 16302 0 16338 25280 4 bl_0_26
port 211 nsew
rlabel metal1 s 16374 0 16410 25280 4 br_0_26
port 213 nsew
rlabel metal1 s 16518 0 16554 25280 4 bl_1_26
port 215 nsew
rlabel metal1 s 16590 0 16626 25280 4 br_1_26
port 217 nsew
rlabel metal1 s 17358 0 17394 25280 4 bl_0_27
port 219 nsew
rlabel metal1 s 17286 0 17322 25280 4 br_0_27
port 221 nsew
rlabel metal1 s 17142 0 17178 25280 4 bl_1_27
port 223 nsew
rlabel metal1 s 17070 0 17106 25280 4 br_1_27
port 225 nsew
rlabel metal1 s 17550 0 17586 25280 4 bl_0_28
port 227 nsew
rlabel metal1 s 17622 0 17658 25280 4 br_0_28
port 229 nsew
rlabel metal1 s 17766 0 17802 25280 4 bl_1_28
port 231 nsew
rlabel metal1 s 17838 0 17874 25280 4 br_1_28
port 233 nsew
rlabel metal1 s 18606 0 18642 25280 4 bl_0_29
port 235 nsew
rlabel metal1 s 18534 0 18570 25280 4 br_0_29
port 237 nsew
rlabel metal1 s 18390 0 18426 25280 4 bl_1_29
port 239 nsew
rlabel metal1 s 18318 0 18354 25280 4 br_1_29
port 241 nsew
rlabel metal1 s 18798 0 18834 25280 4 bl_0_30
port 243 nsew
rlabel metal1 s 18870 0 18906 25280 4 br_0_30
port 245 nsew
rlabel metal1 s 19014 0 19050 25280 4 bl_1_30
port 247 nsew
rlabel metal1 s 19086 0 19122 25280 4 br_1_30
port 249 nsew
rlabel metal1 s 19854 0 19890 25280 4 bl_0_31
port 251 nsew
rlabel metal1 s 19782 0 19818 25280 4 br_0_31
port 253 nsew
rlabel metal1 s 19638 0 19674 25280 4 bl_1_31
port 255 nsew
rlabel metal1 s 19566 0 19602 25280 4 br_1_31
port 257 nsew
rlabel metal2 s 0 323 19968 371 4 wl_0_0
port 259 nsew
rlabel metal2 s 0 103 19968 151 4 wl_1_0
port 261 nsew
rlabel metal2 s 0 419 19968 467 4 wl_0_1
port 263 nsew
rlabel metal2 s 0 639 19968 687 4 wl_1_1
port 265 nsew
rlabel metal2 s 0 1113 19968 1161 4 wl_0_2
port 267 nsew
rlabel metal2 s 0 893 19968 941 4 wl_1_2
port 269 nsew
rlabel metal2 s 0 1209 19968 1257 4 wl_0_3
port 271 nsew
rlabel metal2 s 0 1429 19968 1477 4 wl_1_3
port 273 nsew
rlabel metal2 s 0 1903 19968 1951 4 wl_0_4
port 275 nsew
rlabel metal2 s 0 1683 19968 1731 4 wl_1_4
port 277 nsew
rlabel metal2 s 0 1999 19968 2047 4 wl_0_5
port 279 nsew
rlabel metal2 s 0 2219 19968 2267 4 wl_1_5
port 281 nsew
rlabel metal2 s 0 2693 19968 2741 4 wl_0_6
port 283 nsew
rlabel metal2 s 0 2473 19968 2521 4 wl_1_6
port 285 nsew
rlabel metal2 s 0 2789 19968 2837 4 wl_0_7
port 287 nsew
rlabel metal2 s 0 3009 19968 3057 4 wl_1_7
port 289 nsew
rlabel metal2 s 0 3483 19968 3531 4 wl_0_8
port 291 nsew
rlabel metal2 s 0 3263 19968 3311 4 wl_1_8
port 293 nsew
rlabel metal2 s 0 3579 19968 3627 4 wl_0_9
port 295 nsew
rlabel metal2 s 0 3799 19968 3847 4 wl_1_9
port 297 nsew
rlabel metal2 s 0 4273 19968 4321 4 wl_0_10
port 299 nsew
rlabel metal2 s 0 4053 19968 4101 4 wl_1_10
port 301 nsew
rlabel metal2 s 0 4369 19968 4417 4 wl_0_11
port 303 nsew
rlabel metal2 s 0 4589 19968 4637 4 wl_1_11
port 305 nsew
rlabel metal2 s 0 5063 19968 5111 4 wl_0_12
port 307 nsew
rlabel metal2 s 0 4843 19968 4891 4 wl_1_12
port 309 nsew
rlabel metal2 s 0 5159 19968 5207 4 wl_0_13
port 311 nsew
rlabel metal2 s 0 5379 19968 5427 4 wl_1_13
port 313 nsew
rlabel metal2 s 0 5853 19968 5901 4 wl_0_14
port 315 nsew
rlabel metal2 s 0 5633 19968 5681 4 wl_1_14
port 317 nsew
rlabel metal2 s 0 5949 19968 5997 4 wl_0_15
port 319 nsew
rlabel metal2 s 0 6169 19968 6217 4 wl_1_15
port 321 nsew
rlabel metal2 s 0 6643 19968 6691 4 wl_0_16
port 323 nsew
rlabel metal2 s 0 6423 19968 6471 4 wl_1_16
port 325 nsew
rlabel metal2 s 0 6739 19968 6787 4 wl_0_17
port 327 nsew
rlabel metal2 s 0 6959 19968 7007 4 wl_1_17
port 329 nsew
rlabel metal2 s 0 7433 19968 7481 4 wl_0_18
port 331 nsew
rlabel metal2 s 0 7213 19968 7261 4 wl_1_18
port 333 nsew
rlabel metal2 s 0 7529 19968 7577 4 wl_0_19
port 335 nsew
rlabel metal2 s 0 7749 19968 7797 4 wl_1_19
port 337 nsew
rlabel metal2 s 0 8223 19968 8271 4 wl_0_20
port 339 nsew
rlabel metal2 s 0 8003 19968 8051 4 wl_1_20
port 341 nsew
rlabel metal2 s 0 8319 19968 8367 4 wl_0_21
port 343 nsew
rlabel metal2 s 0 8539 19968 8587 4 wl_1_21
port 345 nsew
rlabel metal2 s 0 9013 19968 9061 4 wl_0_22
port 347 nsew
rlabel metal2 s 0 8793 19968 8841 4 wl_1_22
port 349 nsew
rlabel metal2 s 0 9109 19968 9157 4 wl_0_23
port 351 nsew
rlabel metal2 s 0 9329 19968 9377 4 wl_1_23
port 353 nsew
rlabel metal2 s 0 9803 19968 9851 4 wl_0_24
port 355 nsew
rlabel metal2 s 0 9583 19968 9631 4 wl_1_24
port 357 nsew
rlabel metal2 s 0 9899 19968 9947 4 wl_0_25
port 359 nsew
rlabel metal2 s 0 10119 19968 10167 4 wl_1_25
port 361 nsew
rlabel metal2 s 0 10593 19968 10641 4 wl_0_26
port 363 nsew
rlabel metal2 s 0 10373 19968 10421 4 wl_1_26
port 365 nsew
rlabel metal2 s 0 10689 19968 10737 4 wl_0_27
port 367 nsew
rlabel metal2 s 0 10909 19968 10957 4 wl_1_27
port 369 nsew
rlabel metal2 s 0 11383 19968 11431 4 wl_0_28
port 371 nsew
rlabel metal2 s 0 11163 19968 11211 4 wl_1_28
port 373 nsew
rlabel metal2 s 0 11479 19968 11527 4 wl_0_29
port 375 nsew
rlabel metal2 s 0 11699 19968 11747 4 wl_1_29
port 377 nsew
rlabel metal2 s 0 12173 19968 12221 4 wl_0_30
port 379 nsew
rlabel metal2 s 0 11953 19968 12001 4 wl_1_30
port 381 nsew
rlabel metal2 s 0 12269 19968 12317 4 wl_0_31
port 383 nsew
rlabel metal2 s 0 12489 19968 12537 4 wl_1_31
port 385 nsew
rlabel metal2 s 0 12963 19968 13011 4 wl_0_32
port 387 nsew
rlabel metal2 s 0 12743 19968 12791 4 wl_1_32
port 389 nsew
rlabel metal2 s 0 13059 19968 13107 4 wl_0_33
port 391 nsew
rlabel metal2 s 0 13279 19968 13327 4 wl_1_33
port 393 nsew
rlabel metal2 s 0 13753 19968 13801 4 wl_0_34
port 395 nsew
rlabel metal2 s 0 13533 19968 13581 4 wl_1_34
port 397 nsew
rlabel metal2 s 0 13849 19968 13897 4 wl_0_35
port 399 nsew
rlabel metal2 s 0 14069 19968 14117 4 wl_1_35
port 401 nsew
rlabel metal2 s 0 14543 19968 14591 4 wl_0_36
port 403 nsew
rlabel metal2 s 0 14323 19968 14371 4 wl_1_36
port 405 nsew
rlabel metal2 s 0 14639 19968 14687 4 wl_0_37
port 407 nsew
rlabel metal2 s 0 14859 19968 14907 4 wl_1_37
port 409 nsew
rlabel metal2 s 0 15333 19968 15381 4 wl_0_38
port 411 nsew
rlabel metal2 s 0 15113 19968 15161 4 wl_1_38
port 413 nsew
rlabel metal2 s 0 15429 19968 15477 4 wl_0_39
port 415 nsew
rlabel metal2 s 0 15649 19968 15697 4 wl_1_39
port 417 nsew
rlabel metal2 s 0 16123 19968 16171 4 wl_0_40
port 419 nsew
rlabel metal2 s 0 15903 19968 15951 4 wl_1_40
port 421 nsew
rlabel metal2 s 0 16219 19968 16267 4 wl_0_41
port 423 nsew
rlabel metal2 s 0 16439 19968 16487 4 wl_1_41
port 425 nsew
rlabel metal2 s 0 16913 19968 16961 4 wl_0_42
port 427 nsew
rlabel metal2 s 0 16693 19968 16741 4 wl_1_42
port 429 nsew
rlabel metal2 s 0 17009 19968 17057 4 wl_0_43
port 431 nsew
rlabel metal2 s 0 17229 19968 17277 4 wl_1_43
port 433 nsew
rlabel metal2 s 0 17703 19968 17751 4 wl_0_44
port 435 nsew
rlabel metal2 s 0 17483 19968 17531 4 wl_1_44
port 437 nsew
rlabel metal2 s 0 17799 19968 17847 4 wl_0_45
port 439 nsew
rlabel metal2 s 0 18019 19968 18067 4 wl_1_45
port 441 nsew
rlabel metal2 s 0 18493 19968 18541 4 wl_0_46
port 443 nsew
rlabel metal2 s 0 18273 19968 18321 4 wl_1_46
port 445 nsew
rlabel metal2 s 0 18589 19968 18637 4 wl_0_47
port 447 nsew
rlabel metal2 s 0 18809 19968 18857 4 wl_1_47
port 449 nsew
rlabel metal2 s 0 19283 19968 19331 4 wl_0_48
port 451 nsew
rlabel metal2 s 0 19063 19968 19111 4 wl_1_48
port 453 nsew
rlabel metal2 s 0 19379 19968 19427 4 wl_0_49
port 455 nsew
rlabel metal2 s 0 19599 19968 19647 4 wl_1_49
port 457 nsew
rlabel metal2 s 0 20073 19968 20121 4 wl_0_50
port 459 nsew
rlabel metal2 s 0 19853 19968 19901 4 wl_1_50
port 461 nsew
rlabel metal2 s 0 20169 19968 20217 4 wl_0_51
port 463 nsew
rlabel metal2 s 0 20389 19968 20437 4 wl_1_51
port 465 nsew
rlabel metal2 s 0 20863 19968 20911 4 wl_0_52
port 467 nsew
rlabel metal2 s 0 20643 19968 20691 4 wl_1_52
port 469 nsew
rlabel metal2 s 0 20959 19968 21007 4 wl_0_53
port 471 nsew
rlabel metal2 s 0 21179 19968 21227 4 wl_1_53
port 473 nsew
rlabel metal2 s 0 21653 19968 21701 4 wl_0_54
port 475 nsew
rlabel metal2 s 0 21433 19968 21481 4 wl_1_54
port 477 nsew
rlabel metal2 s 0 21749 19968 21797 4 wl_0_55
port 479 nsew
rlabel metal2 s 0 21969 19968 22017 4 wl_1_55
port 481 nsew
rlabel metal2 s 0 22443 19968 22491 4 wl_0_56
port 483 nsew
rlabel metal2 s 0 22223 19968 22271 4 wl_1_56
port 485 nsew
rlabel metal2 s 0 22539 19968 22587 4 wl_0_57
port 487 nsew
rlabel metal2 s 0 22759 19968 22807 4 wl_1_57
port 489 nsew
rlabel metal2 s 0 23233 19968 23281 4 wl_0_58
port 491 nsew
rlabel metal2 s 0 23013 19968 23061 4 wl_1_58
port 493 nsew
rlabel metal2 s 0 23329 19968 23377 4 wl_0_59
port 495 nsew
rlabel metal2 s 0 23549 19968 23597 4 wl_1_59
port 497 nsew
rlabel metal2 s 0 24023 19968 24071 4 wl_0_60
port 499 nsew
rlabel metal2 s 0 23803 19968 23851 4 wl_1_60
port 501 nsew
rlabel metal2 s 0 24119 19968 24167 4 wl_0_61
port 503 nsew
rlabel metal2 s 0 24339 19968 24387 4 wl_1_61
port 505 nsew
rlabel metal2 s 0 24813 19968 24861 4 wl_0_62
port 507 nsew
rlabel metal2 s 0 24593 19968 24641 4 wl_1_62
port 509 nsew
rlabel metal2 s 0 24909 19968 24957 4 wl_0_63
port 511 nsew
rlabel metal2 s 0 25129 19968 25177 4 wl_1_63
port 513 nsew
rlabel metal1 s 6462 22989 6498 23330 4 vdd
port 515 nsew
rlabel metal1 s 5214 3530 5250 3871 4 vdd
port 515 nsew
rlabel metal1 s 7230 22490 7266 22831 4 vdd
port 515 nsew
rlabel metal1 s 2718 4320 2754 4661 4 vdd
port 515 nsew
rlabel metal1 s 8958 8270 8994 8611 4 vdd
port 515 nsew
rlabel metal1 s 11454 11139 11490 11480 4 vdd
port 515 nsew
rlabel metal1 s 18942 12220 18978 12561 4 vdd
port 515 nsew
rlabel metal1 s 7230 9559 7266 9900 4 vdd
port 515 nsew
rlabel metal1 s 5214 19829 5250 20170 4 vdd
port 515 nsew
rlabel metal1 s 17214 11430 17250 11771 4 vdd
port 515 nsew
rlabel metal1 s 12222 24860 12258 25201 4 vdd
port 515 nsew
rlabel metal1 s 15198 24860 15234 25201 4 vdd
port 515 nsew
rlabel metal1 s 8478 1950 8514 2291 4 vdd
port 515 nsew
rlabel metal1 s 13470 370 13506 711 4 vdd
port 515 nsew
rlabel metal1 s 5982 11139 6018 11480 4 vdd
port 515 nsew
rlabel metal1 s 1470 20619 1506 20960 4 vdd
port 515 nsew
rlabel metal1 s 12222 23280 12258 23621 4 vdd
port 515 nsew
rlabel metal1 s 11454 5900 11490 6241 4 vdd
port 515 nsew
rlabel metal1 s 222 22199 258 22540 4 vdd
port 515 nsew
rlabel metal1 s 11454 14590 11490 14931 4 vdd
port 515 nsew
rlabel metal1 s 17214 11139 17250 11480 4 vdd
port 515 nsew
rlabel metal1 s 11454 8270 11490 8611 4 vdd
port 515 nsew
rlabel metal1 s 11454 8769 11490 9110 4 vdd
port 515 nsew
rlabel metal1 s 14718 13509 14754 13850 4 vdd
port 515 nsew
rlabel metal1 s 15198 1659 15234 2000 4 vdd
port 515 nsew
rlabel metal1 s 14718 20120 14754 20461 4 vdd
port 515 nsew
rlabel metal1 s 11454 22199 11490 22540 4 vdd
port 515 nsew
rlabel metal1 s 8478 4320 8514 4661 4 vdd
port 515 nsew
rlabel metal1 s 2718 16960 2754 17301 4 vdd
port 515 nsew
rlabel metal1 s 8958 1659 8994 2000 4 vdd
port 515 nsew
rlabel metal1 s 6462 20910 6498 21251 4 vdd
port 515 nsew
rlabel metal1 s 11454 6399 11490 6740 4 vdd
port 515 nsew
rlabel metal1 s 15966 17459 16002 17800 4 vdd
port 515 nsew
rlabel metal1 s 5982 20619 6018 20960 4 vdd
port 515 nsew
rlabel metal1 s 18462 1659 18498 2000 4 vdd
port 515 nsew
rlabel metal1 s 8478 11430 8514 11771 4 vdd
port 515 nsew
rlabel metal1 s 12222 14590 12258 14931 4 vdd
port 515 nsew
rlabel metal1 s 17694 8769 17730 9110 4 vdd
port 515 nsew
rlabel metal1 s 3966 20619 4002 20960 4 vdd
port 515 nsew
rlabel metal1 s 13470 23779 13506 24120 4 vdd
port 515 nsew
rlabel metal1 s 13950 8769 13986 9110 4 vdd
port 515 nsew
rlabel metal1 s 7710 9850 7746 10191 4 vdd
port 515 nsew
rlabel metal1 s 12702 22989 12738 23330 4 vdd
port 515 nsew
rlabel metal1 s 5982 5900 6018 6241 4 vdd
port 515 nsew
rlabel metal1 s 19710 16960 19746 17301 4 vdd
port 515 nsew
rlabel metal1 s 18462 11430 18498 11771 4 vdd
port 515 nsew
rlabel metal1 s 2238 23280 2274 23621 4 vdd
port 515 nsew
rlabel metal1 s 14718 6399 14754 6740 4 vdd
port 515 nsew
rlabel metal1 s 16446 22989 16482 23330 4 vdd
port 515 nsew
rlabel metal1 s 10206 10349 10242 10690 4 vdd
port 515 nsew
rlabel metal1 s 15966 12220 16002 12561 4 vdd
port 515 nsew
rlabel metal1 s 10206 7189 10242 7530 4 vdd
port 515 nsew
rlabel metal1 s 11454 21409 11490 21750 4 vdd
port 515 nsew
rlabel metal1 s 18942 3239 18978 3580 4 vdd
port 515 nsew
rlabel metal1 s 990 15879 1026 16220 4 vdd
port 515 nsew
rlabel metal1 s 9726 370 9762 711 4 vdd
port 515 nsew
rlabel metal1 s 18462 15089 18498 15430 4 vdd
port 515 nsew
rlabel metal1 s 9726 12220 9762 12561 4 vdd
port 515 nsew
rlabel metal1 s 222 19330 258 19671 4 vdd
port 515 nsew
rlabel metal1 s 5214 9559 5250 9900 4 vdd
port 515 nsew
rlabel metal1 s 3486 16170 3522 16511 4 vdd
port 515 nsew
rlabel metal1 s 17214 16170 17250 16511 4 vdd
port 515 nsew
rlabel metal1 s 18462 8769 18498 9110 4 vdd
port 515 nsew
rlabel metal1 s 14718 8270 14754 8611 4 vdd
port 515 nsew
rlabel metal1 s 12702 19829 12738 20170 4 vdd
port 515 nsew
rlabel metal1 s 1470 10349 1506 10690 4 vdd
port 515 nsew
rlabel metal1 s 18462 17750 18498 18091 4 vdd
port 515 nsew
rlabel metal1 s 19710 20619 19746 20960 4 vdd
port 515 nsew
rlabel metal1 s 18942 10640 18978 10981 4 vdd
port 515 nsew
rlabel metal1 s 5214 21409 5250 21750 4 vdd
port 515 nsew
rlabel metal1 s 10974 16669 11010 17010 4 vdd
port 515 nsew
rlabel metal1 s 12702 14590 12738 14931 4 vdd
port 515 nsew
rlabel metal1 s 1470 19330 1506 19671 4 vdd
port 515 nsew
rlabel metal1 s 17214 15089 17250 15430 4 vdd
port 515 nsew
rlabel metal1 s 8478 370 8514 711 4 vdd
port 515 nsew
rlabel metal1 s 18942 13800 18978 14141 4 vdd
port 515 nsew
rlabel metal1 s 5982 22490 6018 22831 4 vdd
port 515 nsew
rlabel metal1 s 8478 20120 8514 20461 4 vdd
port 515 nsew
rlabel metal1 s 10974 4320 11010 4661 4 vdd
port 515 nsew
rlabel metal1 s 19710 19330 19746 19671 4 vdd
port 515 nsew
rlabel metal1 s 4734 7189 4770 7530 4 vdd
port 515 nsew
rlabel metal1 s 17214 20120 17250 20461 4 vdd
port 515 nsew
rlabel metal1 s 4734 16669 4770 17010 4 vdd
port 515 nsew
rlabel metal1 s 17694 23779 17730 24120 4 vdd
port 515 nsew
rlabel metal1 s 1470 9060 1506 9401 4 vdd
port 515 nsew
rlabel metal1 s 6462 22199 6498 22540 4 vdd
port 515 nsew
rlabel metal1 s 1470 13509 1506 13850 4 vdd
port 515 nsew
rlabel metal1 s 15198 14299 15234 14640 4 vdd
port 515 nsew
rlabel metal1 s 16446 8769 16482 9110 4 vdd
port 515 nsew
rlabel metal1 s 7230 24569 7266 24910 4 vdd
port 515 nsew
rlabel metal1 s 3966 14299 4002 14640 4 vdd
port 515 nsew
rlabel metal1 s 3966 21409 4002 21750 4 vdd
port 515 nsew
rlabel metal1 s 13950 15879 13986 16220 4 vdd
port 515 nsew
rlabel metal1 s 12702 18540 12738 18881 4 vdd
port 515 nsew
rlabel metal1 s 5214 370 5250 711 4 vdd
port 515 nsew
rlabel metal1 s 1470 23779 1506 24120 4 vdd
port 515 nsew
rlabel metal1 s 13950 9850 13986 10191 4 vdd
port 515 nsew
rlabel metal1 s 12702 15380 12738 15721 4 vdd
port 515 nsew
rlabel metal1 s 15198 7979 15234 8320 4 vdd
port 515 nsew
rlabel metal1 s 3486 11430 3522 11771 4 vdd
port 515 nsew
rlabel metal1 s 3966 16960 4002 17301 4 vdd
port 515 nsew
rlabel metal1 s 15198 19829 15234 20170 4 vdd
port 515 nsew
rlabel metal1 s 222 11430 258 11771 4 vdd
port 515 nsew
rlabel metal1 s 16446 3530 16482 3871 4 vdd
port 515 nsew
rlabel metal1 s 17214 12220 17250 12561 4 vdd
port 515 nsew
rlabel metal1 s 8478 5609 8514 5950 4 vdd
port 515 nsew
rlabel metal1 s 10974 16170 11010 16511 4 vdd
port 515 nsew
rlabel metal1 s 9726 5110 9762 5451 4 vdd
port 515 nsew
rlabel metal1 s 17214 15380 17250 15721 4 vdd
port 515 nsew
rlabel metal1 s 5982 20120 6018 20461 4 vdd
port 515 nsew
rlabel metal1 s 8958 8769 8994 9110 4 vdd
port 515 nsew
rlabel metal1 s 7230 79 7266 420 4 vdd
port 515 nsew
rlabel metal1 s 7230 8769 7266 9110 4 vdd
port 515 nsew
rlabel metal1 s 6462 23779 6498 24120 4 vdd
port 515 nsew
rlabel metal1 s 7710 15879 7746 16220 4 vdd
port 515 nsew
rlabel metal1 s 18462 24860 18498 25201 4 vdd
port 515 nsew
rlabel metal1 s 19710 8270 19746 8611 4 vdd
port 515 nsew
rlabel metal1 s 3966 24860 4002 25201 4 vdd
port 515 nsew
rlabel metal1 s 5214 2740 5250 3081 4 vdd
port 515 nsew
rlabel metal1 s 5214 5609 5250 5950 4 vdd
port 515 nsew
rlabel metal1 s 19710 21700 19746 22041 4 vdd
port 515 nsew
rlabel metal1 s 7230 13509 7266 13850 4 vdd
port 515 nsew
rlabel metal1 s 222 5609 258 5950 4 vdd
port 515 nsew
rlabel metal1 s 3966 8769 4002 9110 4 vdd
port 515 nsew
rlabel metal1 s 19710 5110 19746 5451 4 vdd
port 515 nsew
rlabel metal1 s 14718 2449 14754 2790 4 vdd
port 515 nsew
rlabel metal1 s 7230 20910 7266 21251 4 vdd
port 515 nsew
rlabel metal1 s 12702 17750 12738 18091 4 vdd
port 515 nsew
rlabel metal1 s 6462 24860 6498 25201 4 vdd
port 515 nsew
rlabel metal1 s 12222 19829 12258 20170 4 vdd
port 515 nsew
rlabel metal1 s 10974 370 11010 711 4 vdd
port 515 nsew
rlabel metal1 s 2238 20910 2274 21251 4 vdd
port 515 nsew
rlabel metal1 s 14718 16960 14754 17301 4 vdd
port 515 nsew
rlabel metal1 s 16446 21700 16482 22041 4 vdd
port 515 nsew
rlabel metal1 s 11454 19039 11490 19380 4 vdd
port 515 nsew
rlabel metal1 s 7230 23779 7266 24120 4 vdd
port 515 nsew
rlabel metal1 s 18942 12719 18978 13060 4 vdd
port 515 nsew
rlabel metal1 s 5982 11430 6018 11771 4 vdd
port 515 nsew
rlabel metal1 s 10206 15089 10242 15430 4 vdd
port 515 nsew
rlabel metal1 s 10974 14590 11010 14931 4 vdd
port 515 nsew
rlabel metal1 s 8958 17750 8994 18091 4 vdd
port 515 nsew
rlabel metal1 s 16446 15380 16482 15721 4 vdd
port 515 nsew
rlabel metal1 s 1470 17459 1506 17800 4 vdd
port 515 nsew
rlabel metal1 s 3486 2449 3522 2790 4 vdd
port 515 nsew
rlabel metal1 s 15966 24569 16002 24910 4 vdd
port 515 nsew
rlabel metal1 s 6462 6690 6498 7031 4 vdd
port 515 nsew
rlabel metal1 s 15966 24860 16002 25201 4 vdd
port 515 nsew
rlabel metal1 s 8958 6399 8994 6740 4 vdd
port 515 nsew
rlabel metal1 s 12222 22199 12258 22540 4 vdd
port 515 nsew
rlabel metal1 s 17214 23779 17250 24120 4 vdd
port 515 nsew
rlabel metal1 s 11454 19330 11490 19671 4 vdd
port 515 nsew
rlabel metal1 s 14718 20619 14754 20960 4 vdd
port 515 nsew
rlabel metal1 s 7710 23280 7746 23621 4 vdd
port 515 nsew
rlabel metal1 s 17694 19039 17730 19380 4 vdd
port 515 nsew
rlabel metal1 s 2238 20120 2274 20461 4 vdd
port 515 nsew
rlabel metal1 s 17694 9060 17730 9401 4 vdd
port 515 nsew
rlabel metal1 s 18942 5110 18978 5451 4 vdd
port 515 nsew
rlabel metal1 s 4734 1659 4770 2000 4 vdd
port 515 nsew
rlabel metal1 s 18942 13010 18978 13351 4 vdd
port 515 nsew
rlabel metal1 s 19710 2449 19746 2790 4 vdd
port 515 nsew
rlabel metal1 s 4734 13509 4770 13850 4 vdd
port 515 nsew
rlabel metal1 s 17694 6399 17730 6740 4 vdd
port 515 nsew
rlabel metal1 s 5214 6690 5250 7031 4 vdd
port 515 nsew
rlabel metal1 s 222 24860 258 25201 4 vdd
port 515 nsew
rlabel metal1 s 19710 21409 19746 21750 4 vdd
port 515 nsew
rlabel metal1 s 5982 5609 6018 5950 4 vdd
port 515 nsew
rlabel metal1 s 6462 7979 6498 8320 4 vdd
port 515 nsew
rlabel metal1 s 11454 13010 11490 13351 4 vdd
port 515 nsew
rlabel metal1 s 14718 13800 14754 14141 4 vdd
port 515 nsew
rlabel metal1 s 13950 9559 13986 9900 4 vdd
port 515 nsew
rlabel metal1 s 9726 10349 9762 10690 4 vdd
port 515 nsew
rlabel metal1 s 17694 11139 17730 11480 4 vdd
port 515 nsew
rlabel metal1 s 15966 3239 16002 3580 4 vdd
port 515 nsew
rlabel metal1 s 12702 869 12738 1210 4 vdd
port 515 nsew
rlabel metal1 s 10974 13509 11010 13850 4 vdd
port 515 nsew
rlabel metal1 s 16446 22490 16482 22831 4 vdd
port 515 nsew
rlabel metal1 s 222 370 258 711 4 vdd
port 515 nsew
rlabel metal1 s 9726 9559 9762 9900 4 vdd
port 515 nsew
rlabel metal1 s 18462 6690 18498 7031 4 vdd
port 515 nsew
rlabel metal1 s 10206 6399 10242 6740 4 vdd
port 515 nsew
rlabel metal1 s 2718 9060 2754 9401 4 vdd
port 515 nsew
rlabel metal1 s 9726 15380 9762 15721 4 vdd
port 515 nsew
rlabel metal1 s 19710 3239 19746 3580 4 vdd
port 515 nsew
rlabel metal1 s 7710 9060 7746 9401 4 vdd
port 515 nsew
rlabel metal1 s 6462 10349 6498 10690 4 vdd
port 515 nsew
rlabel metal1 s 13950 16669 13986 17010 4 vdd
port 515 nsew
rlabel metal1 s 19710 15380 19746 15721 4 vdd
port 515 nsew
rlabel metal1 s 12702 1659 12738 2000 4 vdd
port 515 nsew
rlabel metal1 s 14718 21409 14754 21750 4 vdd
port 515 nsew
rlabel metal1 s 17214 19039 17250 19380 4 vdd
port 515 nsew
rlabel metal1 s 19710 370 19746 711 4 vdd
port 515 nsew
rlabel metal1 s 17214 19829 17250 20170 4 vdd
port 515 nsew
rlabel metal1 s 17214 7480 17250 7821 4 vdd
port 515 nsew
rlabel metal1 s 12702 13800 12738 14141 4 vdd
port 515 nsew
rlabel metal1 s 15966 9850 16002 10191 4 vdd
port 515 nsew
rlabel metal1 s 9726 11929 9762 12270 4 vdd
port 515 nsew
rlabel metal1 s 17214 5609 17250 5950 4 vdd
port 515 nsew
rlabel metal1 s 10206 869 10242 1210 4 vdd
port 515 nsew
rlabel metal1 s 15198 17459 15234 17800 4 vdd
port 515 nsew
rlabel metal1 s 5982 3530 6018 3871 4 vdd
port 515 nsew
rlabel metal1 s 6462 10640 6498 10981 4 vdd
port 515 nsew
rlabel metal1 s 13950 24070 13986 24411 4 vdd
port 515 nsew
rlabel metal1 s 7230 15089 7266 15430 4 vdd
port 515 nsew
rlabel metal1 s 11454 14299 11490 14640 4 vdd
port 515 nsew
rlabel metal1 s 8958 15879 8994 16220 4 vdd
port 515 nsew
rlabel metal1 s 6462 16960 6498 17301 4 vdd
port 515 nsew
rlabel metal1 s 2238 23779 2274 24120 4 vdd
port 515 nsew
rlabel metal1 s 18942 24569 18978 24910 4 vdd
port 515 nsew
rlabel metal1 s 3966 869 4002 1210 4 vdd
port 515 nsew
rlabel metal1 s 5214 18540 5250 18881 4 vdd
port 515 nsew
rlabel metal1 s 8478 21700 8514 22041 4 vdd
port 515 nsew
rlabel metal1 s 17694 22989 17730 23330 4 vdd
port 515 nsew
rlabel metal1 s 8958 18540 8994 18881 4 vdd
port 515 nsew
rlabel metal1 s 4734 6690 4770 7031 4 vdd
port 515 nsew
rlabel metal1 s 2238 6690 2274 7031 4 vdd
port 515 nsew
rlabel metal1 s 9726 13010 9762 13351 4 vdd
port 515 nsew
rlabel metal1 s 18942 16669 18978 17010 4 vdd
port 515 nsew
rlabel metal1 s 8958 1950 8994 2291 4 vdd
port 515 nsew
rlabel metal1 s 17694 15089 17730 15430 4 vdd
port 515 nsew
rlabel metal1 s 12222 11139 12258 11480 4 vdd
port 515 nsew
rlabel metal1 s 12222 3239 12258 3580 4 vdd
port 515 nsew
rlabel metal1 s 15966 11430 16002 11771 4 vdd
port 515 nsew
rlabel metal1 s 10974 79 11010 420 4 vdd
port 515 nsew
rlabel metal1 s 3486 869 3522 1210 4 vdd
port 515 nsew
rlabel metal1 s 12702 12220 12738 12561 4 vdd
port 515 nsew
rlabel metal1 s 13470 6690 13506 7031 4 vdd
port 515 nsew
rlabel metal1 s 6462 869 6498 1210 4 vdd
port 515 nsew
rlabel metal1 s 11454 12719 11490 13060 4 vdd
port 515 nsew
rlabel metal1 s 2718 21409 2754 21750 4 vdd
port 515 nsew
rlabel metal1 s 3966 13800 4002 14141 4 vdd
port 515 nsew
rlabel metal1 s 9726 19829 9762 20170 4 vdd
port 515 nsew
rlabel metal1 s 2718 13800 2754 14141 4 vdd
port 515 nsew
rlabel metal1 s 5214 8769 5250 9110 4 vdd
port 515 nsew
rlabel metal1 s 4734 9850 4770 10191 4 vdd
port 515 nsew
rlabel metal1 s 222 1160 258 1501 4 vdd
port 515 nsew
rlabel metal1 s 8478 21409 8514 21750 4 vdd
port 515 nsew
rlabel metal1 s 18942 7189 18978 7530 4 vdd
port 515 nsew
rlabel metal1 s 7710 15380 7746 15721 4 vdd
port 515 nsew
rlabel metal1 s 3966 13010 4002 13351 4 vdd
port 515 nsew
rlabel metal1 s 17694 14590 17730 14931 4 vdd
port 515 nsew
rlabel metal1 s 13950 11929 13986 12270 4 vdd
port 515 nsew
rlabel metal1 s 6462 20619 6498 20960 4 vdd
port 515 nsew
rlabel metal1 s 13950 21409 13986 21750 4 vdd
port 515 nsew
rlabel metal1 s 8958 6690 8994 7031 4 vdd
port 515 nsew
rlabel metal1 s 17694 20910 17730 21251 4 vdd
port 515 nsew
rlabel metal1 s 8478 10640 8514 10981 4 vdd
port 515 nsew
rlabel metal1 s 5982 12220 6018 12561 4 vdd
port 515 nsew
rlabel metal1 s 4734 16170 4770 16511 4 vdd
port 515 nsew
rlabel metal1 s 18462 24569 18498 24910 4 vdd
port 515 nsew
rlabel metal1 s 5982 16170 6018 16511 4 vdd
port 515 nsew
rlabel metal1 s 13470 19829 13506 20170 4 vdd
port 515 nsew
rlabel metal1 s 10206 22989 10242 23330 4 vdd
port 515 nsew
rlabel metal1 s 16446 869 16482 1210 4 vdd
port 515 nsew
rlabel metal1 s 12222 10640 12258 10981 4 vdd
port 515 nsew
rlabel metal1 s 7230 4029 7266 4370 4 vdd
port 515 nsew
rlabel metal1 s 1470 7979 1506 8320 4 vdd
port 515 nsew
rlabel metal1 s 9726 79 9762 420 4 vdd
port 515 nsew
rlabel metal1 s 14718 18249 14754 18590 4 vdd
port 515 nsew
rlabel metal1 s 15198 5110 15234 5451 4 vdd
port 515 nsew
rlabel metal1 s 14718 18540 14754 18881 4 vdd
port 515 nsew
rlabel metal1 s 4734 9559 4770 9900 4 vdd
port 515 nsew
rlabel metal1 s 4734 3239 4770 3580 4 vdd
port 515 nsew
rlabel metal1 s 2238 17750 2274 18091 4 vdd
port 515 nsew
rlabel metal1 s 12222 12220 12258 12561 4 vdd
port 515 nsew
rlabel metal1 s 13470 14590 13506 14931 4 vdd
port 515 nsew
rlabel metal1 s 4734 14590 4770 14931 4 vdd
port 515 nsew
rlabel metal1 s 222 22989 258 23330 4 vdd
port 515 nsew
rlabel metal1 s 11454 22490 11490 22831 4 vdd
port 515 nsew
rlabel metal1 s 10206 3239 10242 3580 4 vdd
port 515 nsew
rlabel metal1 s 11454 24569 11490 24910 4 vdd
port 515 nsew
rlabel metal1 s 18462 2449 18498 2790 4 vdd
port 515 nsew
rlabel metal1 s 4734 4819 4770 5160 4 vdd
port 515 nsew
rlabel metal1 s 18462 3239 18498 3580 4 vdd
port 515 nsew
rlabel metal1 s 5982 16960 6018 17301 4 vdd
port 515 nsew
rlabel metal1 s 17694 21409 17730 21750 4 vdd
port 515 nsew
rlabel metal1 s 15966 16170 16002 16511 4 vdd
port 515 nsew
rlabel metal1 s 12222 16170 12258 16511 4 vdd
port 515 nsew
rlabel metal1 s 3486 22199 3522 22540 4 vdd
port 515 nsew
rlabel metal1 s 4734 21700 4770 22041 4 vdd
port 515 nsew
rlabel metal1 s 12702 21409 12738 21750 4 vdd
port 515 nsew
rlabel metal1 s 7230 23280 7266 23621 4 vdd
port 515 nsew
rlabel metal1 s 19710 20910 19746 21251 4 vdd
port 515 nsew
rlabel metal1 s 5982 17750 6018 18091 4 vdd
port 515 nsew
rlabel metal1 s 7710 23779 7746 24120 4 vdd
port 515 nsew
rlabel metal1 s 17694 5110 17730 5451 4 vdd
port 515 nsew
rlabel metal1 s 990 16960 1026 17301 4 vdd
port 515 nsew
rlabel metal1 s 4734 11929 4770 12270 4 vdd
port 515 nsew
rlabel metal1 s 18942 869 18978 1210 4 vdd
port 515 nsew
rlabel metal1 s 5982 1160 6018 1501 4 vdd
port 515 nsew
rlabel metal1 s 3966 10640 4002 10981 4 vdd
port 515 nsew
rlabel metal1 s 990 18540 1026 18881 4 vdd
port 515 nsew
rlabel metal1 s 17214 24070 17250 24411 4 vdd
port 515 nsew
rlabel metal1 s 18942 4029 18978 4370 4 vdd
port 515 nsew
rlabel metal1 s 10206 4320 10242 4661 4 vdd
port 515 nsew
rlabel metal1 s 13950 20120 13986 20461 4 vdd
port 515 nsew
rlabel metal1 s 16446 16960 16482 17301 4 vdd
port 515 nsew
rlabel metal1 s 18462 10349 18498 10690 4 vdd
port 515 nsew
rlabel metal1 s 15966 17750 16002 18091 4 vdd
port 515 nsew
rlabel metal1 s 5214 79 5250 420 4 vdd
port 515 nsew
rlabel metal1 s 5982 20910 6018 21251 4 vdd
port 515 nsew
rlabel metal1 s 990 7480 1026 7821 4 vdd
port 515 nsew
rlabel metal1 s 8958 16170 8994 16511 4 vdd
port 515 nsew
rlabel metal1 s 3966 18249 4002 18590 4 vdd
port 515 nsew
rlabel metal1 s 9726 2449 9762 2790 4 vdd
port 515 nsew
rlabel metal1 s 3486 1160 3522 1501 4 vdd
port 515 nsew
rlabel metal1 s 16446 1160 16482 1501 4 vdd
port 515 nsew
rlabel metal1 s 7230 19330 7266 19671 4 vdd
port 515 nsew
rlabel metal1 s 13470 10640 13506 10981 4 vdd
port 515 nsew
rlabel metal1 s 990 7979 1026 8320 4 vdd
port 515 nsew
rlabel metal1 s 11454 5609 11490 5950 4 vdd
port 515 nsew
rlabel metal1 s 16446 4029 16482 4370 4 vdd
port 515 nsew
rlabel metal1 s 10974 17750 11010 18091 4 vdd
port 515 nsew
rlabel metal1 s 10974 6399 11010 6740 4 vdd
port 515 nsew
rlabel metal1 s 18462 20120 18498 20461 4 vdd
port 515 nsew
rlabel metal1 s 12222 17750 12258 18091 4 vdd
port 515 nsew
rlabel metal1 s 6462 9850 6498 10191 4 vdd
port 515 nsew
rlabel metal1 s 3486 8270 3522 8611 4 vdd
port 515 nsew
rlabel metal1 s 18462 7979 18498 8320 4 vdd
port 515 nsew
rlabel metal1 s 18942 15089 18978 15430 4 vdd
port 515 nsew
rlabel metal1 s 18462 19330 18498 19671 4 vdd
port 515 nsew
rlabel metal1 s 13950 10640 13986 10981 4 vdd
port 515 nsew
rlabel metal1 s 12222 3530 12258 3871 4 vdd
port 515 nsew
rlabel metal1 s 16446 13509 16482 13850 4 vdd
port 515 nsew
rlabel metal1 s 7710 21700 7746 22041 4 vdd
port 515 nsew
rlabel metal1 s 2238 7979 2274 8320 4 vdd
port 515 nsew
rlabel metal1 s 15198 22199 15234 22540 4 vdd
port 515 nsew
rlabel metal1 s 17214 13509 17250 13850 4 vdd
port 515 nsew
rlabel metal1 s 5214 1659 5250 2000 4 vdd
port 515 nsew
rlabel metal1 s 1470 13010 1506 13351 4 vdd
port 515 nsew
rlabel metal1 s 13470 11139 13506 11480 4 vdd
port 515 nsew
rlabel metal1 s 12222 20120 12258 20461 4 vdd
port 515 nsew
rlabel metal1 s 8478 16669 8514 17010 4 vdd
port 515 nsew
rlabel metal1 s 5982 12719 6018 13060 4 vdd
port 515 nsew
rlabel metal1 s 5982 22199 6018 22540 4 vdd
port 515 nsew
rlabel metal1 s 990 869 1026 1210 4 vdd
port 515 nsew
rlabel metal1 s 2718 9559 2754 9900 4 vdd
port 515 nsew
rlabel metal1 s 11454 6690 11490 7031 4 vdd
port 515 nsew
rlabel metal1 s 17694 79 17730 420 4 vdd
port 515 nsew
rlabel metal1 s 18462 13800 18498 14141 4 vdd
port 515 nsew
rlabel metal1 s 17694 7189 17730 7530 4 vdd
port 515 nsew
rlabel metal1 s 2718 16669 2754 17010 4 vdd
port 515 nsew
rlabel metal1 s 18942 6399 18978 6740 4 vdd
port 515 nsew
rlabel metal1 s 7230 22989 7266 23330 4 vdd
port 515 nsew
rlabel metal1 s 11454 18249 11490 18590 4 vdd
port 515 nsew
rlabel metal1 s 7230 5900 7266 6241 4 vdd
port 515 nsew
rlabel metal1 s 15198 16669 15234 17010 4 vdd
port 515 nsew
rlabel metal1 s 16446 5900 16482 6241 4 vdd
port 515 nsew
rlabel metal1 s 222 10349 258 10690 4 vdd
port 515 nsew
rlabel metal1 s 10206 15380 10242 15721 4 vdd
port 515 nsew
rlabel metal1 s 4734 4320 4770 4661 4 vdd
port 515 nsew
rlabel metal1 s 16446 16170 16482 16511 4 vdd
port 515 nsew
rlabel metal1 s 10206 15879 10242 16220 4 vdd
port 515 nsew
rlabel metal1 s 10206 19330 10242 19671 4 vdd
port 515 nsew
rlabel metal1 s 13470 12220 13506 12561 4 vdd
port 515 nsew
rlabel metal1 s 5982 7979 6018 8320 4 vdd
port 515 nsew
rlabel metal1 s 15966 16960 16002 17301 4 vdd
port 515 nsew
rlabel metal1 s 222 11929 258 12270 4 vdd
port 515 nsew
rlabel metal1 s 3966 15089 4002 15430 4 vdd
port 515 nsew
rlabel metal1 s 11454 11929 11490 12270 4 vdd
port 515 nsew
rlabel metal1 s 15198 5609 15234 5950 4 vdd
port 515 nsew
rlabel metal1 s 13470 3530 13506 3871 4 vdd
port 515 nsew
rlabel metal1 s 17694 3530 17730 3871 4 vdd
port 515 nsew
rlabel metal1 s 15198 7189 15234 7530 4 vdd
port 515 nsew
rlabel metal1 s 2238 14299 2274 14640 4 vdd
port 515 nsew
rlabel metal1 s 16446 19330 16482 19671 4 vdd
port 515 nsew
rlabel metal1 s 222 2449 258 2790 4 vdd
port 515 nsew
rlabel metal1 s 16446 4320 16482 4661 4 vdd
port 515 nsew
rlabel metal1 s 2238 24070 2274 24411 4 vdd
port 515 nsew
rlabel metal1 s 7710 3530 7746 3871 4 vdd
port 515 nsew
rlabel metal1 s 16446 79 16482 420 4 vdd
port 515 nsew
rlabel metal1 s 8478 14299 8514 14640 4 vdd
port 515 nsew
rlabel metal1 s 13470 22989 13506 23330 4 vdd
port 515 nsew
rlabel metal1 s 1470 18249 1506 18590 4 vdd
port 515 nsew
rlabel metal1 s 19710 5609 19746 5950 4 vdd
port 515 nsew
rlabel metal1 s 8958 7979 8994 8320 4 vdd
port 515 nsew
rlabel metal1 s 19710 10349 19746 10690 4 vdd
port 515 nsew
rlabel metal1 s 3966 10349 4002 10690 4 vdd
port 515 nsew
rlabel metal1 s 11454 18540 11490 18881 4 vdd
port 515 nsew
rlabel metal1 s 16446 10640 16482 10981 4 vdd
port 515 nsew
rlabel metal1 s 2718 2449 2754 2790 4 vdd
port 515 nsew
rlabel metal1 s 3966 23779 4002 24120 4 vdd
port 515 nsew
rlabel metal1 s 10206 1659 10242 2000 4 vdd
port 515 nsew
rlabel metal1 s 6462 18249 6498 18590 4 vdd
port 515 nsew
rlabel metal1 s 7230 11430 7266 11771 4 vdd
port 515 nsew
rlabel metal1 s 7230 11929 7266 12270 4 vdd
port 515 nsew
rlabel metal1 s 10206 11430 10242 11771 4 vdd
port 515 nsew
rlabel metal1 s 18942 79 18978 420 4 vdd
port 515 nsew
rlabel metal1 s 990 22199 1026 22540 4 vdd
port 515 nsew
rlabel metal1 s 7710 16170 7746 16511 4 vdd
port 515 nsew
rlabel metal1 s 12222 869 12258 1210 4 vdd
port 515 nsew
rlabel metal1 s 13470 13800 13506 14141 4 vdd
port 515 nsew
rlabel metal1 s 18942 18249 18978 18590 4 vdd
port 515 nsew
rlabel metal1 s 18462 24070 18498 24411 4 vdd
port 515 nsew
rlabel metal1 s 222 19039 258 19380 4 vdd
port 515 nsew
rlabel metal1 s 12702 11929 12738 12270 4 vdd
port 515 nsew
rlabel metal1 s 7230 5110 7266 5451 4 vdd
port 515 nsew
rlabel metal1 s 6462 1659 6498 2000 4 vdd
port 515 nsew
rlabel metal1 s 14718 12220 14754 12561 4 vdd
port 515 nsew
rlabel metal1 s 2238 5900 2274 6241 4 vdd
port 515 nsew
rlabel metal1 s 18462 19039 18498 19380 4 vdd
port 515 nsew
rlabel metal1 s 3486 5900 3522 6241 4 vdd
port 515 nsew
rlabel metal1 s 15198 12719 15234 13060 4 vdd
port 515 nsew
rlabel metal1 s 12222 13010 12258 13351 4 vdd
port 515 nsew
rlabel metal1 s 14718 24569 14754 24910 4 vdd
port 515 nsew
rlabel metal1 s 8478 6399 8514 6740 4 vdd
port 515 nsew
rlabel metal1 s 2718 4029 2754 4370 4 vdd
port 515 nsew
rlabel metal1 s 17694 16960 17730 17301 4 vdd
port 515 nsew
rlabel metal1 s 13950 24569 13986 24910 4 vdd
port 515 nsew
rlabel metal1 s 5214 16960 5250 17301 4 vdd
port 515 nsew
rlabel metal1 s 9726 18249 9762 18590 4 vdd
port 515 nsew
rlabel metal1 s 5982 8769 6018 9110 4 vdd
port 515 nsew
rlabel metal1 s 12702 22490 12738 22831 4 vdd
port 515 nsew
rlabel metal1 s 18942 11139 18978 11480 4 vdd
port 515 nsew
rlabel metal1 s 18462 7480 18498 7821 4 vdd
port 515 nsew
rlabel metal1 s 2718 9850 2754 10191 4 vdd
port 515 nsew
rlabel metal1 s 14718 10640 14754 10981 4 vdd
port 515 nsew
rlabel metal1 s 9726 3530 9762 3871 4 vdd
port 515 nsew
rlabel metal1 s 10206 14590 10242 14931 4 vdd
port 515 nsew
rlabel metal1 s 15198 79 15234 420 4 vdd
port 515 nsew
rlabel metal1 s 12702 12719 12738 13060 4 vdd
port 515 nsew
rlabel metal1 s 7710 2449 7746 2790 4 vdd
port 515 nsew
rlabel metal1 s 2718 10640 2754 10981 4 vdd
port 515 nsew
rlabel metal1 s 7710 11929 7746 12270 4 vdd
port 515 nsew
rlabel metal1 s 8958 2740 8994 3081 4 vdd
port 515 nsew
rlabel metal1 s 10206 9850 10242 10191 4 vdd
port 515 nsew
rlabel metal1 s 8478 24070 8514 24411 4 vdd
port 515 nsew
rlabel metal1 s 6462 7189 6498 7530 4 vdd
port 515 nsew
rlabel metal1 s 7230 12719 7266 13060 4 vdd
port 515 nsew
rlabel metal1 s 11454 24070 11490 24411 4 vdd
port 515 nsew
rlabel metal1 s 10974 10349 11010 10690 4 vdd
port 515 nsew
rlabel metal1 s 5214 5110 5250 5451 4 vdd
port 515 nsew
rlabel metal1 s 13950 79 13986 420 4 vdd
port 515 nsew
rlabel metal1 s 11454 4320 11490 4661 4 vdd
port 515 nsew
rlabel metal1 s 10974 2449 11010 2790 4 vdd
port 515 nsew
rlabel metal1 s 12222 21700 12258 22041 4 vdd
port 515 nsew
rlabel metal1 s 15966 14590 16002 14931 4 vdd
port 515 nsew
rlabel metal1 s 222 13800 258 14141 4 vdd
port 515 nsew
rlabel metal1 s 1470 20120 1506 20461 4 vdd
port 515 nsew
rlabel metal1 s 13950 15380 13986 15721 4 vdd
port 515 nsew
rlabel metal1 s 4734 15879 4770 16220 4 vdd
port 515 nsew
rlabel metal1 s 7230 9060 7266 9401 4 vdd
port 515 nsew
rlabel metal1 s 12702 8769 12738 9110 4 vdd
port 515 nsew
rlabel metal1 s 2718 20120 2754 20461 4 vdd
port 515 nsew
rlabel metal1 s 12222 5609 12258 5950 4 vdd
port 515 nsew
rlabel metal1 s 5982 1950 6018 2291 4 vdd
port 515 nsew
rlabel metal1 s 18942 370 18978 711 4 vdd
port 515 nsew
rlabel metal1 s 13950 13010 13986 13351 4 vdd
port 515 nsew
rlabel metal1 s 13470 11430 13506 11771 4 vdd
port 515 nsew
rlabel metal1 s 15198 3530 15234 3871 4 vdd
port 515 nsew
rlabel metal1 s 7710 18249 7746 18590 4 vdd
port 515 nsew
rlabel metal1 s 15966 22199 16002 22540 4 vdd
port 515 nsew
rlabel metal1 s 8958 3530 8994 3871 4 vdd
port 515 nsew
rlabel metal1 s 12222 11430 12258 11771 4 vdd
port 515 nsew
rlabel metal1 s 12702 4029 12738 4370 4 vdd
port 515 nsew
rlabel metal1 s 15198 9850 15234 10191 4 vdd
port 515 nsew
rlabel metal1 s 18462 14299 18498 14640 4 vdd
port 515 nsew
rlabel metal1 s 17694 9850 17730 10191 4 vdd
port 515 nsew
rlabel metal1 s 10206 4029 10242 4370 4 vdd
port 515 nsew
rlabel metal1 s 10206 19039 10242 19380 4 vdd
port 515 nsew
rlabel metal1 s 16446 7189 16482 7530 4 vdd
port 515 nsew
rlabel metal1 s 14718 5110 14754 5451 4 vdd
port 515 nsew
rlabel metal1 s 3966 5609 4002 5950 4 vdd
port 515 nsew
rlabel metal1 s 13470 20910 13506 21251 4 vdd
port 515 nsew
rlabel metal1 s 15966 19330 16002 19671 4 vdd
port 515 nsew
rlabel metal1 s 10206 6690 10242 7031 4 vdd
port 515 nsew
rlabel metal1 s 19710 16669 19746 17010 4 vdd
port 515 nsew
rlabel metal1 s 990 15089 1026 15430 4 vdd
port 515 nsew
rlabel metal1 s 8958 24569 8994 24910 4 vdd
port 515 nsew
rlabel metal1 s 4734 22490 4770 22831 4 vdd
port 515 nsew
rlabel metal1 s 18462 16170 18498 16511 4 vdd
port 515 nsew
rlabel metal1 s 5982 14590 6018 14931 4 vdd
port 515 nsew
rlabel metal1 s 3486 15879 3522 16220 4 vdd
port 515 nsew
rlabel metal1 s 2718 370 2754 711 4 vdd
port 515 nsew
rlabel metal1 s 12222 8270 12258 8611 4 vdd
port 515 nsew
rlabel metal1 s 5982 9850 6018 10191 4 vdd
port 515 nsew
rlabel metal1 s 15198 18249 15234 18590 4 vdd
port 515 nsew
rlabel metal1 s 222 4029 258 4370 4 vdd
port 515 nsew
rlabel metal1 s 16446 2449 16482 2790 4 vdd
port 515 nsew
rlabel metal1 s 15966 21700 16002 22041 4 vdd
port 515 nsew
rlabel metal1 s 8478 869 8514 1210 4 vdd
port 515 nsew
rlabel metal1 s 5214 14590 5250 14931 4 vdd
port 515 nsew
rlabel metal1 s 5982 19039 6018 19380 4 vdd
port 515 nsew
rlabel metal1 s 12222 20910 12258 21251 4 vdd
port 515 nsew
rlabel metal1 s 5982 23779 6018 24120 4 vdd
port 515 nsew
rlabel metal1 s 15966 19039 16002 19380 4 vdd
port 515 nsew
rlabel metal1 s 990 17459 1026 17800 4 vdd
port 515 nsew
rlabel metal1 s 10974 19039 11010 19380 4 vdd
port 515 nsew
rlabel metal1 s 3486 4320 3522 4661 4 vdd
port 515 nsew
rlabel metal1 s 13470 10349 13506 10690 4 vdd
port 515 nsew
rlabel metal1 s 7710 22490 7746 22831 4 vdd
port 515 nsew
rlabel metal1 s 222 1659 258 2000 4 vdd
port 515 nsew
rlabel metal1 s 16446 9559 16482 9900 4 vdd
port 515 nsew
rlabel metal1 s 6462 4320 6498 4661 4 vdd
port 515 nsew
rlabel metal1 s 11454 370 11490 711 4 vdd
port 515 nsew
rlabel metal1 s 8958 79 8994 420 4 vdd
port 515 nsew
rlabel metal1 s 12222 16960 12258 17301 4 vdd
port 515 nsew
rlabel metal1 s 3966 22989 4002 23330 4 vdd
port 515 nsew
rlabel metal1 s 9726 16669 9762 17010 4 vdd
port 515 nsew
rlabel metal1 s 7710 4819 7746 5160 4 vdd
port 515 nsew
rlabel metal1 s 13950 21700 13986 22041 4 vdd
port 515 nsew
rlabel metal1 s 18462 11929 18498 12270 4 vdd
port 515 nsew
rlabel metal1 s 18942 23779 18978 24120 4 vdd
port 515 nsew
rlabel metal1 s 17214 4029 17250 4370 4 vdd
port 515 nsew
rlabel metal1 s 10974 4819 11010 5160 4 vdd
port 515 nsew
rlabel metal1 s 3486 79 3522 420 4 vdd
port 515 nsew
rlabel metal1 s 5214 20619 5250 20960 4 vdd
port 515 nsew
rlabel metal1 s 18942 1160 18978 1501 4 vdd
port 515 nsew
rlabel metal1 s 11454 23280 11490 23621 4 vdd
port 515 nsew
rlabel metal1 s 16446 8270 16482 8611 4 vdd
port 515 nsew
rlabel metal1 s 13950 7189 13986 7530 4 vdd
port 515 nsew
rlabel metal1 s 990 79 1026 420 4 vdd
port 515 nsew
rlabel metal1 s 2718 23280 2754 23621 4 vdd
port 515 nsew
rlabel metal1 s 2718 24569 2754 24910 4 vdd
port 515 nsew
rlabel metal1 s 8478 6690 8514 7031 4 vdd
port 515 nsew
rlabel metal1 s 15966 20619 16002 20960 4 vdd
port 515 nsew
rlabel metal1 s 18462 79 18498 420 4 vdd
port 515 nsew
rlabel metal1 s 8478 4819 8514 5160 4 vdd
port 515 nsew
rlabel metal1 s 9726 22989 9762 23330 4 vdd
port 515 nsew
rlabel metal1 s 4734 79 4770 420 4 vdd
port 515 nsew
rlabel metal1 s 3966 9559 4002 9900 4 vdd
port 515 nsew
rlabel metal1 s 15966 12719 16002 13060 4 vdd
port 515 nsew
rlabel metal1 s 10974 11139 11010 11480 4 vdd
port 515 nsew
rlabel metal1 s 7230 2449 7266 2790 4 vdd
port 515 nsew
rlabel metal1 s 18462 7189 18498 7530 4 vdd
port 515 nsew
rlabel metal1 s 7230 24860 7266 25201 4 vdd
port 515 nsew
rlabel metal1 s 1470 15089 1506 15430 4 vdd
port 515 nsew
rlabel metal1 s 5982 5110 6018 5451 4 vdd
port 515 nsew
rlabel metal1 s 222 22490 258 22831 4 vdd
port 515 nsew
rlabel metal1 s 12222 13509 12258 13850 4 vdd
port 515 nsew
rlabel metal1 s 990 1160 1026 1501 4 vdd
port 515 nsew
rlabel metal1 s 6462 11929 6498 12270 4 vdd
port 515 nsew
rlabel metal1 s 990 4029 1026 4370 4 vdd
port 515 nsew
rlabel metal1 s 3486 7979 3522 8320 4 vdd
port 515 nsew
rlabel metal1 s 17694 9559 17730 9900 4 vdd
port 515 nsew
rlabel metal1 s 6462 370 6498 711 4 vdd
port 515 nsew
rlabel metal1 s 12702 15879 12738 16220 4 vdd
port 515 nsew
rlabel metal1 s 15198 370 15234 711 4 vdd
port 515 nsew
rlabel metal1 s 12222 2449 12258 2790 4 vdd
port 515 nsew
rlabel metal1 s 12702 22199 12738 22540 4 vdd
port 515 nsew
rlabel metal1 s 7230 10349 7266 10690 4 vdd
port 515 nsew
rlabel metal1 s 2718 24070 2754 24411 4 vdd
port 515 nsew
rlabel metal1 s 15966 13509 16002 13850 4 vdd
port 515 nsew
rlabel metal1 s 12702 20619 12738 20960 4 vdd
port 515 nsew
rlabel metal1 s 13470 869 13506 1210 4 vdd
port 515 nsew
rlabel metal1 s 990 23779 1026 24120 4 vdd
port 515 nsew
rlabel metal1 s 10974 8270 11010 8611 4 vdd
port 515 nsew
rlabel metal1 s 11454 13800 11490 14141 4 vdd
port 515 nsew
rlabel metal1 s 3486 18540 3522 18881 4 vdd
port 515 nsew
rlabel metal1 s 7230 19039 7266 19380 4 vdd
port 515 nsew
rlabel metal1 s 19710 22490 19746 22831 4 vdd
port 515 nsew
rlabel metal1 s 3966 7189 4002 7530 4 vdd
port 515 nsew
rlabel metal1 s 17214 3530 17250 3871 4 vdd
port 515 nsew
rlabel metal1 s 4734 19829 4770 20170 4 vdd
port 515 nsew
rlabel metal1 s 13950 16170 13986 16511 4 vdd
port 515 nsew
rlabel metal1 s 6462 11139 6498 11480 4 vdd
port 515 nsew
rlabel metal1 s 3486 11139 3522 11480 4 vdd
port 515 nsew
rlabel metal1 s 2238 15089 2274 15430 4 vdd
port 515 nsew
rlabel metal1 s 13470 4029 13506 4370 4 vdd
port 515 nsew
rlabel metal1 s 3966 8270 4002 8611 4 vdd
port 515 nsew
rlabel metal1 s 13950 20619 13986 20960 4 vdd
port 515 nsew
rlabel metal1 s 7710 19330 7746 19671 4 vdd
port 515 nsew
rlabel metal1 s 11454 20619 11490 20960 4 vdd
port 515 nsew
rlabel metal1 s 13950 12220 13986 12561 4 vdd
port 515 nsew
rlabel metal1 s 990 18249 1026 18590 4 vdd
port 515 nsew
rlabel metal1 s 3966 9060 4002 9401 4 vdd
port 515 nsew
rlabel metal1 s 7710 20120 7746 20461 4 vdd
port 515 nsew
rlabel metal1 s 4734 18249 4770 18590 4 vdd
port 515 nsew
rlabel metal1 s 6462 3530 6498 3871 4 vdd
port 515 nsew
rlabel metal1 s 13950 20910 13986 21251 4 vdd
port 515 nsew
rlabel metal1 s 7710 6399 7746 6740 4 vdd
port 515 nsew
rlabel metal1 s 8478 23280 8514 23621 4 vdd
port 515 nsew
rlabel metal1 s 990 6690 1026 7031 4 vdd
port 515 nsew
rlabel metal1 s 10974 11929 11010 12270 4 vdd
port 515 nsew
rlabel metal1 s 12222 370 12258 711 4 vdd
port 515 nsew
rlabel metal1 s 15198 15089 15234 15430 4 vdd
port 515 nsew
rlabel metal1 s 10974 19330 11010 19671 4 vdd
port 515 nsew
rlabel metal1 s 11454 24860 11490 25201 4 vdd
port 515 nsew
rlabel metal1 s 19710 10640 19746 10981 4 vdd
port 515 nsew
rlabel metal1 s 2718 5900 2754 6241 4 vdd
port 515 nsew
rlabel metal1 s 1470 24070 1506 24411 4 vdd
port 515 nsew
rlabel metal1 s 2718 18540 2754 18881 4 vdd
port 515 nsew
rlabel metal1 s 8958 19829 8994 20170 4 vdd
port 515 nsew
rlabel metal1 s 8478 5110 8514 5451 4 vdd
port 515 nsew
rlabel metal1 s 2718 22490 2754 22831 4 vdd
port 515 nsew
rlabel metal1 s 1470 14299 1506 14640 4 vdd
port 515 nsew
rlabel metal1 s 10206 5110 10242 5451 4 vdd
port 515 nsew
rlabel metal1 s 16446 14590 16482 14931 4 vdd
port 515 nsew
rlabel metal1 s 10206 24860 10242 25201 4 vdd
port 515 nsew
rlabel metal1 s 7230 13010 7266 13351 4 vdd
port 515 nsew
rlabel metal1 s 7710 16960 7746 17301 4 vdd
port 515 nsew
rlabel metal1 s 18462 13509 18498 13850 4 vdd
port 515 nsew
rlabel metal1 s 18942 19039 18978 19380 4 vdd
port 515 nsew
rlabel metal1 s 8478 13800 8514 14141 4 vdd
port 515 nsew
rlabel metal1 s 5214 7480 5250 7821 4 vdd
port 515 nsew
rlabel metal1 s 7710 10349 7746 10690 4 vdd
port 515 nsew
rlabel metal1 s 222 12719 258 13060 4 vdd
port 515 nsew
rlabel metal1 s 18462 4320 18498 4661 4 vdd
port 515 nsew
rlabel metal1 s 15966 3530 16002 3871 4 vdd
port 515 nsew
rlabel metal1 s 4734 12719 4770 13060 4 vdd
port 515 nsew
rlabel metal1 s 1470 9850 1506 10191 4 vdd
port 515 nsew
rlabel metal1 s 5214 11929 5250 12270 4 vdd
port 515 nsew
rlabel metal1 s 990 19330 1026 19671 4 vdd
port 515 nsew
rlabel metal1 s 17694 19829 17730 20170 4 vdd
port 515 nsew
rlabel metal1 s 3486 6690 3522 7031 4 vdd
port 515 nsew
rlabel metal1 s 15966 8769 16002 9110 4 vdd
port 515 nsew
rlabel metal1 s 12702 4819 12738 5160 4 vdd
port 515 nsew
rlabel metal1 s 5214 18249 5250 18590 4 vdd
port 515 nsew
rlabel metal1 s 5982 16669 6018 17010 4 vdd
port 515 nsew
rlabel metal1 s 990 8270 1026 8611 4 vdd
port 515 nsew
rlabel metal1 s 15198 4320 15234 4661 4 vdd
port 515 nsew
rlabel metal1 s 7710 11430 7746 11771 4 vdd
port 515 nsew
rlabel metal1 s 10974 5609 11010 5950 4 vdd
port 515 nsew
rlabel metal1 s 15198 16960 15234 17301 4 vdd
port 515 nsew
rlabel metal1 s 2718 19330 2754 19671 4 vdd
port 515 nsew
rlabel metal1 s 5214 4029 5250 4370 4 vdd
port 515 nsew
rlabel metal1 s 12222 2740 12258 3081 4 vdd
port 515 nsew
rlabel metal1 s 8958 14590 8994 14931 4 vdd
port 515 nsew
rlabel metal1 s 1470 14590 1506 14931 4 vdd
port 515 nsew
rlabel metal1 s 8958 19330 8994 19671 4 vdd
port 515 nsew
rlabel metal1 s 15198 16170 15234 16511 4 vdd
port 515 nsew
rlabel metal1 s 17214 22989 17250 23330 4 vdd
port 515 nsew
rlabel metal1 s 990 24860 1026 25201 4 vdd
port 515 nsew
rlabel metal1 s 1470 8270 1506 8611 4 vdd
port 515 nsew
rlabel metal1 s 18462 15380 18498 15721 4 vdd
port 515 nsew
rlabel metal1 s 12702 17459 12738 17800 4 vdd
port 515 nsew
rlabel metal1 s 7230 18540 7266 18881 4 vdd
port 515 nsew
rlabel metal1 s 222 2740 258 3081 4 vdd
port 515 nsew
rlabel metal1 s 1470 22199 1506 22540 4 vdd
port 515 nsew
rlabel metal1 s 10206 23280 10242 23621 4 vdd
port 515 nsew
rlabel metal1 s 222 9850 258 10191 4 vdd
port 515 nsew
rlabel metal1 s 2718 22199 2754 22540 4 vdd
port 515 nsew
rlabel metal1 s 18942 5609 18978 5950 4 vdd
port 515 nsew
rlabel metal1 s 13470 7979 13506 8320 4 vdd
port 515 nsew
rlabel metal1 s 18462 16669 18498 17010 4 vdd
port 515 nsew
rlabel metal1 s 10206 22490 10242 22831 4 vdd
port 515 nsew
rlabel metal1 s 8478 18249 8514 18590 4 vdd
port 515 nsew
rlabel metal1 s 18462 9850 18498 10191 4 vdd
port 515 nsew
rlabel metal1 s 9726 17750 9762 18091 4 vdd
port 515 nsew
rlabel metal1 s 10974 21700 11010 22041 4 vdd
port 515 nsew
rlabel metal1 s 10974 9850 11010 10191 4 vdd
port 515 nsew
rlabel metal1 s 11454 7480 11490 7821 4 vdd
port 515 nsew
rlabel metal1 s 12702 1950 12738 2291 4 vdd
port 515 nsew
rlabel metal1 s 18942 17459 18978 17800 4 vdd
port 515 nsew
rlabel metal1 s 18942 7979 18978 8320 4 vdd
port 515 nsew
rlabel metal1 s 13950 3239 13986 3580 4 vdd
port 515 nsew
rlabel metal1 s 8958 3239 8994 3580 4 vdd
port 515 nsew
rlabel metal1 s 19710 7480 19746 7821 4 vdd
port 515 nsew
rlabel metal1 s 3966 4320 4002 4661 4 vdd
port 515 nsew
rlabel metal1 s 17694 4819 17730 5160 4 vdd
port 515 nsew
rlabel metal1 s 13470 5609 13506 5950 4 vdd
port 515 nsew
rlabel metal1 s 15966 4320 16002 4661 4 vdd
port 515 nsew
rlabel metal1 s 7710 10640 7746 10981 4 vdd
port 515 nsew
rlabel metal1 s 12702 13010 12738 13351 4 vdd
port 515 nsew
rlabel metal1 s 17694 15380 17730 15721 4 vdd
port 515 nsew
rlabel metal1 s 15966 1659 16002 2000 4 vdd
port 515 nsew
rlabel metal1 s 4734 11139 4770 11480 4 vdd
port 515 nsew
rlabel metal1 s 9726 21700 9762 22041 4 vdd
port 515 nsew
rlabel metal1 s 1470 6690 1506 7031 4 vdd
port 515 nsew
rlabel metal1 s 3966 1659 4002 2000 4 vdd
port 515 nsew
rlabel metal1 s 5982 21409 6018 21750 4 vdd
port 515 nsew
rlabel metal1 s 11454 10640 11490 10981 4 vdd
port 515 nsew
rlabel metal1 s 12222 4819 12258 5160 4 vdd
port 515 nsew
rlabel metal1 s 8958 19039 8994 19380 4 vdd
port 515 nsew
rlabel metal1 s 16446 19039 16482 19380 4 vdd
port 515 nsew
rlabel metal1 s 10206 8270 10242 8611 4 vdd
port 515 nsew
rlabel metal1 s 5214 9060 5250 9401 4 vdd
port 515 nsew
rlabel metal1 s 10206 13800 10242 14141 4 vdd
port 515 nsew
rlabel metal1 s 3486 19829 3522 20170 4 vdd
port 515 nsew
rlabel metal1 s 5982 24569 6018 24910 4 vdd
port 515 nsew
rlabel metal1 s 3486 10349 3522 10690 4 vdd
port 515 nsew
rlabel metal1 s 10206 2449 10242 2790 4 vdd
port 515 nsew
rlabel metal1 s 12222 1950 12258 2291 4 vdd
port 515 nsew
rlabel metal1 s 10974 12719 11010 13060 4 vdd
port 515 nsew
rlabel metal1 s 2238 9060 2274 9401 4 vdd
port 515 nsew
rlabel metal1 s 4734 3530 4770 3871 4 vdd
port 515 nsew
rlabel metal1 s 15198 15380 15234 15721 4 vdd
port 515 nsew
rlabel metal1 s 13470 12719 13506 13060 4 vdd
port 515 nsew
rlabel metal1 s 5214 15089 5250 15430 4 vdd
port 515 nsew
rlabel metal1 s 8958 20120 8994 20461 4 vdd
port 515 nsew
rlabel metal1 s 9726 14299 9762 14640 4 vdd
port 515 nsew
rlabel metal1 s 222 20619 258 20960 4 vdd
port 515 nsew
rlabel metal1 s 10974 3530 11010 3871 4 vdd
port 515 nsew
rlabel metal1 s 8478 7979 8514 8320 4 vdd
port 515 nsew
rlabel metal1 s 2238 6399 2274 6740 4 vdd
port 515 nsew
rlabel metal1 s 8958 10640 8994 10981 4 vdd
port 515 nsew
rlabel metal1 s 16446 9850 16482 10191 4 vdd
port 515 nsew
rlabel metal1 s 3966 11929 4002 12270 4 vdd
port 515 nsew
rlabel metal1 s 3486 17750 3522 18091 4 vdd
port 515 nsew
rlabel metal1 s 10974 24070 11010 24411 4 vdd
port 515 nsew
rlabel metal1 s 6462 14299 6498 14640 4 vdd
port 515 nsew
rlabel metal1 s 7230 9850 7266 10191 4 vdd
port 515 nsew
rlabel metal1 s 9726 12719 9762 13060 4 vdd
port 515 nsew
rlabel metal1 s 10974 20910 11010 21251 4 vdd
port 515 nsew
rlabel metal1 s 4734 2449 4770 2790 4 vdd
port 515 nsew
rlabel metal1 s 10974 19829 11010 20170 4 vdd
port 515 nsew
rlabel metal1 s 11454 15380 11490 15721 4 vdd
port 515 nsew
rlabel metal1 s 3486 20619 3522 20960 4 vdd
port 515 nsew
rlabel metal1 s 2718 6690 2754 7031 4 vdd
port 515 nsew
rlabel metal1 s 14718 22490 14754 22831 4 vdd
port 515 nsew
rlabel metal1 s 8478 15380 8514 15721 4 vdd
port 515 nsew
rlabel metal1 s 12222 20619 12258 20960 4 vdd
port 515 nsew
rlabel metal1 s 17214 7189 17250 7530 4 vdd
port 515 nsew
rlabel metal1 s 18942 24860 18978 25201 4 vdd
port 515 nsew
rlabel metal1 s 990 5609 1026 5950 4 vdd
port 515 nsew
rlabel metal1 s 1470 869 1506 1210 4 vdd
port 515 nsew
rlabel metal1 s 2718 14590 2754 14931 4 vdd
port 515 nsew
rlabel metal1 s 3966 17750 4002 18091 4 vdd
port 515 nsew
rlabel metal1 s 2718 14299 2754 14640 4 vdd
port 515 nsew
rlabel metal1 s 2238 16960 2274 17301 4 vdd
port 515 nsew
rlabel metal1 s 13950 19829 13986 20170 4 vdd
port 515 nsew
rlabel metal1 s 18462 4819 18498 5160 4 vdd
port 515 nsew
rlabel metal1 s 222 7979 258 8320 4 vdd
port 515 nsew
rlabel metal1 s 14718 11139 14754 11480 4 vdd
port 515 nsew
rlabel metal1 s 3486 9060 3522 9401 4 vdd
port 515 nsew
rlabel metal1 s 7230 22199 7266 22540 4 vdd
port 515 nsew
rlabel metal1 s 13950 19039 13986 19380 4 vdd
port 515 nsew
rlabel metal1 s 8478 4029 8514 4370 4 vdd
port 515 nsew
rlabel metal1 s 13470 23280 13506 23621 4 vdd
port 515 nsew
rlabel metal1 s 11454 11430 11490 11771 4 vdd
port 515 nsew
rlabel metal1 s 7230 5609 7266 5950 4 vdd
port 515 nsew
rlabel metal1 s 14718 9850 14754 10191 4 vdd
port 515 nsew
rlabel metal1 s 15966 4819 16002 5160 4 vdd
port 515 nsew
rlabel metal1 s 3486 21700 3522 22041 4 vdd
port 515 nsew
rlabel metal1 s 10206 18540 10242 18881 4 vdd
port 515 nsew
rlabel metal1 s 13950 2740 13986 3081 4 vdd
port 515 nsew
rlabel metal1 s 16446 12220 16482 12561 4 vdd
port 515 nsew
rlabel metal1 s 4734 12220 4770 12561 4 vdd
port 515 nsew
rlabel metal1 s 17694 869 17730 1210 4 vdd
port 515 nsew
rlabel metal1 s 6462 8270 6498 8611 4 vdd
port 515 nsew
rlabel metal1 s 15966 1950 16002 2291 4 vdd
port 515 nsew
rlabel metal1 s 15198 13800 15234 14141 4 vdd
port 515 nsew
rlabel metal1 s 18942 13509 18978 13850 4 vdd
port 515 nsew
rlabel metal1 s 2718 1160 2754 1501 4 vdd
port 515 nsew
rlabel metal1 s 990 9850 1026 10191 4 vdd
port 515 nsew
rlabel metal1 s 17694 7480 17730 7821 4 vdd
port 515 nsew
rlabel metal1 s 18462 22490 18498 22831 4 vdd
port 515 nsew
rlabel metal1 s 990 14299 1026 14640 4 vdd
port 515 nsew
rlabel metal1 s 2238 16669 2274 17010 4 vdd
port 515 nsew
rlabel metal1 s 18942 20619 18978 20960 4 vdd
port 515 nsew
rlabel metal1 s 5982 15089 6018 15430 4 vdd
port 515 nsew
rlabel metal1 s 2238 9559 2274 9900 4 vdd
port 515 nsew
rlabel metal1 s 18942 2740 18978 3081 4 vdd
port 515 nsew
rlabel metal1 s 18462 22199 18498 22540 4 vdd
port 515 nsew
rlabel metal1 s 14718 24070 14754 24411 4 vdd
port 515 nsew
rlabel metal1 s 13950 17459 13986 17800 4 vdd
port 515 nsew
rlabel metal1 s 3966 19330 4002 19671 4 vdd
port 515 nsew
rlabel metal1 s 15966 2740 16002 3081 4 vdd
port 515 nsew
rlabel metal1 s 15966 20120 16002 20461 4 vdd
port 515 nsew
rlabel metal1 s 8478 7480 8514 7821 4 vdd
port 515 nsew
rlabel metal1 s 16446 5609 16482 5950 4 vdd
port 515 nsew
rlabel metal1 s 3966 1160 4002 1501 4 vdd
port 515 nsew
rlabel metal1 s 10206 22199 10242 22540 4 vdd
port 515 nsew
rlabel metal1 s 11454 4819 11490 5160 4 vdd
port 515 nsew
rlabel metal1 s 990 16669 1026 17010 4 vdd
port 515 nsew
rlabel metal1 s 9726 13509 9762 13850 4 vdd
port 515 nsew
rlabel metal1 s 8958 5900 8994 6241 4 vdd
port 515 nsew
rlabel metal1 s 3486 24070 3522 24411 4 vdd
port 515 nsew
rlabel metal1 s 2718 8270 2754 8611 4 vdd
port 515 nsew
rlabel metal1 s 2238 3239 2274 3580 4 vdd
port 515 nsew
rlabel metal1 s 12702 16170 12738 16511 4 vdd
port 515 nsew
rlabel metal1 s 10206 21700 10242 22041 4 vdd
port 515 nsew
rlabel metal1 s 12222 14299 12258 14640 4 vdd
port 515 nsew
rlabel metal1 s 13470 9559 13506 9900 4 vdd
port 515 nsew
rlabel metal1 s 8478 17750 8514 18091 4 vdd
port 515 nsew
rlabel metal1 s 12702 4320 12738 4661 4 vdd
port 515 nsew
rlabel metal1 s 8958 11929 8994 12270 4 vdd
port 515 nsew
rlabel metal1 s 2718 24860 2754 25201 4 vdd
port 515 nsew
rlabel metal1 s 6462 4029 6498 4370 4 vdd
port 515 nsew
rlabel metal1 s 3486 3239 3522 3580 4 vdd
port 515 nsew
rlabel metal1 s 990 14590 1026 14931 4 vdd
port 515 nsew
rlabel metal1 s 6462 1160 6498 1501 4 vdd
port 515 nsew
rlabel metal1 s 19710 24569 19746 24910 4 vdd
port 515 nsew
rlabel metal1 s 12702 11139 12738 11480 4 vdd
port 515 nsew
rlabel metal1 s 1470 2740 1506 3081 4 vdd
port 515 nsew
rlabel metal1 s 10206 370 10242 711 4 vdd
port 515 nsew
rlabel metal1 s 6462 19039 6498 19380 4 vdd
port 515 nsew
rlabel metal1 s 17214 21700 17250 22041 4 vdd
port 515 nsew
rlabel metal1 s 15198 20120 15234 20461 4 vdd
port 515 nsew
rlabel metal1 s 12702 3239 12738 3580 4 vdd
port 515 nsew
rlabel metal1 s 1470 5900 1506 6241 4 vdd
port 515 nsew
rlabel metal1 s 14718 15089 14754 15430 4 vdd
port 515 nsew
rlabel metal1 s 17214 13800 17250 14141 4 vdd
port 515 nsew
rlabel metal1 s 10206 9559 10242 9900 4 vdd
port 515 nsew
rlabel metal1 s 19710 22199 19746 22540 4 vdd
port 515 nsew
rlabel metal1 s 16446 23280 16482 23621 4 vdd
port 515 nsew
rlabel metal1 s 8478 19330 8514 19671 4 vdd
port 515 nsew
rlabel metal1 s 12702 9850 12738 10191 4 vdd
port 515 nsew
rlabel metal1 s 5214 22989 5250 23330 4 vdd
port 515 nsew
rlabel metal1 s 12702 7480 12738 7821 4 vdd
port 515 nsew
rlabel metal1 s 9726 23779 9762 24120 4 vdd
port 515 nsew
rlabel metal1 s 6462 22490 6498 22831 4 vdd
port 515 nsew
rlabel metal1 s 5982 79 6018 420 4 vdd
port 515 nsew
rlabel metal1 s 10974 10640 11010 10981 4 vdd
port 515 nsew
rlabel metal1 s 15966 16669 16002 17010 4 vdd
port 515 nsew
rlabel metal1 s 10974 20120 11010 20461 4 vdd
port 515 nsew
rlabel metal1 s 1470 79 1506 420 4 vdd
port 515 nsew
rlabel metal1 s 5214 1950 5250 2291 4 vdd
port 515 nsew
rlabel metal1 s 13470 5110 13506 5451 4 vdd
port 515 nsew
rlabel metal1 s 18942 19330 18978 19671 4 vdd
port 515 nsew
rlabel metal1 s 18462 6399 18498 6740 4 vdd
port 515 nsew
rlabel metal1 s 12702 2449 12738 2790 4 vdd
port 515 nsew
rlabel metal1 s 222 9060 258 9401 4 vdd
port 515 nsew
rlabel metal1 s 990 10349 1026 10690 4 vdd
port 515 nsew
rlabel metal1 s 13950 1659 13986 2000 4 vdd
port 515 nsew
rlabel metal1 s 15198 869 15234 1210 4 vdd
port 515 nsew
rlabel metal1 s 8958 24070 8994 24411 4 vdd
port 515 nsew
rlabel metal1 s 5214 14299 5250 14640 4 vdd
port 515 nsew
rlabel metal1 s 14718 7189 14754 7530 4 vdd
port 515 nsew
rlabel metal1 s 15966 10349 16002 10690 4 vdd
port 515 nsew
rlabel metal1 s 2238 13509 2274 13850 4 vdd
port 515 nsew
rlabel metal1 s 17214 11929 17250 12270 4 vdd
port 515 nsew
rlabel metal1 s 222 21700 258 22041 4 vdd
port 515 nsew
rlabel metal1 s 18942 1950 18978 2291 4 vdd
port 515 nsew
rlabel metal1 s 11454 1160 11490 1501 4 vdd
port 515 nsew
rlabel metal1 s 10206 7480 10242 7821 4 vdd
port 515 nsew
rlabel metal1 s 15198 10349 15234 10690 4 vdd
port 515 nsew
rlabel metal1 s 13470 19039 13506 19380 4 vdd
port 515 nsew
rlabel metal1 s 9726 20120 9762 20461 4 vdd
port 515 nsew
rlabel metal1 s 19710 4819 19746 5160 4 vdd
port 515 nsew
rlabel metal1 s 4734 1950 4770 2291 4 vdd
port 515 nsew
rlabel metal1 s 9726 7189 9762 7530 4 vdd
port 515 nsew
rlabel metal1 s 18462 11139 18498 11480 4 vdd
port 515 nsew
rlabel metal1 s 4734 10349 4770 10690 4 vdd
port 515 nsew
rlabel metal1 s 2238 13800 2274 14141 4 vdd
port 515 nsew
rlabel metal1 s 19710 14590 19746 14931 4 vdd
port 515 nsew
rlabel metal1 s 12702 5110 12738 5451 4 vdd
port 515 nsew
rlabel metal1 s 5982 18249 6018 18590 4 vdd
port 515 nsew
rlabel metal1 s 17214 23280 17250 23621 4 vdd
port 515 nsew
rlabel metal1 s 11454 3530 11490 3871 4 vdd
port 515 nsew
rlabel metal1 s 17214 7979 17250 8320 4 vdd
port 515 nsew
rlabel metal1 s 7710 5609 7746 5950 4 vdd
port 515 nsew
rlabel metal1 s 7710 5900 7746 6241 4 vdd
port 515 nsew
rlabel metal1 s 17694 16170 17730 16511 4 vdd
port 515 nsew
rlabel metal1 s 9726 24860 9762 25201 4 vdd
port 515 nsew
rlabel metal1 s 2238 1160 2274 1501 4 vdd
port 515 nsew
rlabel metal1 s 18462 9559 18498 9900 4 vdd
port 515 nsew
rlabel metal1 s 11454 7979 11490 8320 4 vdd
port 515 nsew
rlabel metal1 s 10974 12220 11010 12561 4 vdd
port 515 nsew
rlabel metal1 s 15198 17750 15234 18091 4 vdd
port 515 nsew
rlabel metal1 s 9726 22490 9762 22831 4 vdd
port 515 nsew
rlabel metal1 s 15966 23779 16002 24120 4 vdd
port 515 nsew
rlabel metal1 s 8478 9850 8514 10191 4 vdd
port 515 nsew
rlabel metal1 s 2718 12719 2754 13060 4 vdd
port 515 nsew
rlabel metal1 s 5214 11139 5250 11480 4 vdd
port 515 nsew
rlabel metal1 s 17694 5900 17730 6241 4 vdd
port 515 nsew
rlabel metal1 s 990 3239 1026 3580 4 vdd
port 515 nsew
rlabel metal1 s 13470 21409 13506 21750 4 vdd
port 515 nsew
rlabel metal1 s 9726 15089 9762 15430 4 vdd
port 515 nsew
rlabel metal1 s 6462 21409 6498 21750 4 vdd
port 515 nsew
rlabel metal1 s 7230 14299 7266 14640 4 vdd
port 515 nsew
rlabel metal1 s 10974 22989 11010 23330 4 vdd
port 515 nsew
rlabel metal1 s 990 12220 1026 12561 4 vdd
port 515 nsew
rlabel metal1 s 12222 24569 12258 24910 4 vdd
port 515 nsew
rlabel metal1 s 8958 10349 8994 10690 4 vdd
port 515 nsew
rlabel metal1 s 15966 8270 16002 8611 4 vdd
port 515 nsew
rlabel metal1 s 7710 2740 7746 3081 4 vdd
port 515 nsew
rlabel metal1 s 222 6690 258 7031 4 vdd
port 515 nsew
rlabel metal1 s 5982 2449 6018 2790 4 vdd
port 515 nsew
rlabel metal1 s 2238 21409 2274 21750 4 vdd
port 515 nsew
rlabel metal1 s 14718 15879 14754 16220 4 vdd
port 515 nsew
rlabel metal1 s 13950 10349 13986 10690 4 vdd
port 515 nsew
rlabel metal1 s 8958 15380 8994 15721 4 vdd
port 515 nsew
rlabel metal1 s 6462 17459 6498 17800 4 vdd
port 515 nsew
rlabel metal1 s 11454 17459 11490 17800 4 vdd
port 515 nsew
rlabel metal1 s 13950 22989 13986 23330 4 vdd
port 515 nsew
rlabel metal1 s 5214 13800 5250 14141 4 vdd
port 515 nsew
rlabel metal1 s 17694 11430 17730 11771 4 vdd
port 515 nsew
rlabel metal1 s 12702 19039 12738 19380 4 vdd
port 515 nsew
rlabel metal1 s 990 7189 1026 7530 4 vdd
port 515 nsew
rlabel metal1 s 1470 370 1506 711 4 vdd
port 515 nsew
rlabel metal1 s 14718 22989 14754 23330 4 vdd
port 515 nsew
rlabel metal1 s 7230 15380 7266 15721 4 vdd
port 515 nsew
rlabel metal1 s 3966 11139 4002 11480 4 vdd
port 515 nsew
rlabel metal1 s 13470 7480 13506 7821 4 vdd
port 515 nsew
rlabel metal1 s 2238 4320 2274 4661 4 vdd
port 515 nsew
rlabel metal1 s 18462 5609 18498 5950 4 vdd
port 515 nsew
rlabel metal1 s 3966 4819 4002 5160 4 vdd
port 515 nsew
rlabel metal1 s 10974 6690 11010 7031 4 vdd
port 515 nsew
rlabel metal1 s 15198 12220 15234 12561 4 vdd
port 515 nsew
rlabel metal1 s 15966 5110 16002 5451 4 vdd
port 515 nsew
rlabel metal1 s 10974 23779 11010 24120 4 vdd
port 515 nsew
rlabel metal1 s 15198 20910 15234 21251 4 vdd
port 515 nsew
rlabel metal1 s 19710 19829 19746 20170 4 vdd
port 515 nsew
rlabel metal1 s 12222 6690 12258 7031 4 vdd
port 515 nsew
rlabel metal1 s 12222 24070 12258 24411 4 vdd
port 515 nsew
rlabel metal1 s 19710 6399 19746 6740 4 vdd
port 515 nsew
rlabel metal1 s 8958 7189 8994 7530 4 vdd
port 515 nsew
rlabel metal1 s 2238 370 2274 711 4 vdd
port 515 nsew
rlabel metal1 s 17694 6690 17730 7031 4 vdd
port 515 nsew
rlabel metal1 s 18462 9060 18498 9401 4 vdd
port 515 nsew
rlabel metal1 s 9726 4029 9762 4370 4 vdd
port 515 nsew
rlabel metal1 s 8478 22199 8514 22540 4 vdd
port 515 nsew
rlabel metal1 s 3486 13800 3522 14141 4 vdd
port 515 nsew
rlabel metal1 s 3966 24070 4002 24411 4 vdd
port 515 nsew
rlabel metal1 s 5214 869 5250 1210 4 vdd
port 515 nsew
rlabel metal1 s 2238 11139 2274 11480 4 vdd
port 515 nsew
rlabel metal1 s 5214 1160 5250 1501 4 vdd
port 515 nsew
rlabel metal1 s 13470 6399 13506 6740 4 vdd
port 515 nsew
rlabel metal1 s 11454 869 11490 1210 4 vdd
port 515 nsew
rlabel metal1 s 8478 24860 8514 25201 4 vdd
port 515 nsew
rlabel metal1 s 16446 1950 16482 2291 4 vdd
port 515 nsew
rlabel metal1 s 10206 8769 10242 9110 4 vdd
port 515 nsew
rlabel metal1 s 990 20910 1026 21251 4 vdd
port 515 nsew
rlabel metal1 s 15966 15380 16002 15721 4 vdd
port 515 nsew
rlabel metal1 s 3486 23779 3522 24120 4 vdd
port 515 nsew
rlabel metal1 s 6462 19330 6498 19671 4 vdd
port 515 nsew
rlabel metal1 s 4734 17750 4770 18091 4 vdd
port 515 nsew
rlabel metal1 s 17214 3239 17250 3580 4 vdd
port 515 nsew
rlabel metal1 s 3486 6399 3522 6740 4 vdd
port 515 nsew
rlabel metal1 s 15966 9060 16002 9401 4 vdd
port 515 nsew
rlabel metal1 s 3966 20910 4002 21251 4 vdd
port 515 nsew
rlabel metal1 s 222 15879 258 16220 4 vdd
port 515 nsew
rlabel metal1 s 1470 18540 1506 18881 4 vdd
port 515 nsew
rlabel metal1 s 16446 2740 16482 3081 4 vdd
port 515 nsew
rlabel metal1 s 19710 17459 19746 17800 4 vdd
port 515 nsew
rlabel metal1 s 10206 1160 10242 1501 4 vdd
port 515 nsew
rlabel metal1 s 10206 14299 10242 14640 4 vdd
port 515 nsew
rlabel metal1 s 8478 16170 8514 16511 4 vdd
port 515 nsew
rlabel metal1 s 18462 23779 18498 24120 4 vdd
port 515 nsew
rlabel metal1 s 990 2449 1026 2790 4 vdd
port 515 nsew
rlabel metal1 s 990 20120 1026 20461 4 vdd
port 515 nsew
rlabel metal1 s 13950 7979 13986 8320 4 vdd
port 515 nsew
rlabel metal1 s 3486 9850 3522 10191 4 vdd
port 515 nsew
rlabel metal1 s 14718 22199 14754 22540 4 vdd
port 515 nsew
rlabel metal1 s 8958 4819 8994 5160 4 vdd
port 515 nsew
rlabel metal1 s 19710 11929 19746 12270 4 vdd
port 515 nsew
rlabel metal1 s 15966 370 16002 711 4 vdd
port 515 nsew
rlabel metal1 s 13470 4819 13506 5160 4 vdd
port 515 nsew
rlabel metal1 s 13950 7480 13986 7821 4 vdd
port 515 nsew
rlabel metal1 s 4734 24569 4770 24910 4 vdd
port 515 nsew
rlabel metal1 s 3966 16170 4002 16511 4 vdd
port 515 nsew
rlabel metal1 s 7230 11139 7266 11480 4 vdd
port 515 nsew
rlabel metal1 s 17214 21409 17250 21750 4 vdd
port 515 nsew
rlabel metal1 s 222 4320 258 4661 4 vdd
port 515 nsew
rlabel metal1 s 2238 24860 2274 25201 4 vdd
port 515 nsew
rlabel metal1 s 8478 13509 8514 13850 4 vdd
port 515 nsew
rlabel metal1 s 1470 16960 1506 17301 4 vdd
port 515 nsew
rlabel metal1 s 7230 17750 7266 18091 4 vdd
port 515 nsew
rlabel metal1 s 17214 5900 17250 6241 4 vdd
port 515 nsew
rlabel metal1 s 1470 5110 1506 5451 4 vdd
port 515 nsew
rlabel metal1 s 10974 13800 11010 14141 4 vdd
port 515 nsew
rlabel metal1 s 9726 23280 9762 23621 4 vdd
port 515 nsew
rlabel metal1 s 11454 9060 11490 9401 4 vdd
port 515 nsew
rlabel metal1 s 3966 24569 4002 24910 4 vdd
port 515 nsew
rlabel metal1 s 7230 18249 7266 18590 4 vdd
port 515 nsew
rlabel metal1 s 10974 13010 11010 13351 4 vdd
port 515 nsew
rlabel metal1 s 15966 18540 16002 18881 4 vdd
port 515 nsew
rlabel metal1 s 15966 79 16002 420 4 vdd
port 515 nsew
rlabel metal1 s 18942 22989 18978 23330 4 vdd
port 515 nsew
rlabel metal1 s 10974 17459 11010 17800 4 vdd
port 515 nsew
rlabel metal1 s 222 12220 258 12561 4 vdd
port 515 nsew
rlabel metal1 s 7710 20910 7746 21251 4 vdd
port 515 nsew
rlabel metal1 s 13470 15089 13506 15430 4 vdd
port 515 nsew
rlabel metal1 s 12222 10349 12258 10690 4 vdd
port 515 nsew
rlabel metal1 s 15198 13010 15234 13351 4 vdd
port 515 nsew
rlabel metal1 s 10974 16960 11010 17301 4 vdd
port 515 nsew
rlabel metal1 s 18942 14299 18978 14640 4 vdd
port 515 nsew
rlabel metal1 s 1470 4320 1506 4661 4 vdd
port 515 nsew
rlabel metal1 s 13950 1160 13986 1501 4 vdd
port 515 nsew
rlabel metal1 s 5982 11929 6018 12270 4 vdd
port 515 nsew
rlabel metal1 s 990 9060 1026 9401 4 vdd
port 515 nsew
rlabel metal1 s 18942 7480 18978 7821 4 vdd
port 515 nsew
rlabel metal1 s 17694 18249 17730 18590 4 vdd
port 515 nsew
rlabel metal1 s 18462 13010 18498 13351 4 vdd
port 515 nsew
rlabel metal1 s 3486 24860 3522 25201 4 vdd
port 515 nsew
rlabel metal1 s 11454 16960 11490 17301 4 vdd
port 515 nsew
rlabel metal1 s 14718 19039 14754 19380 4 vdd
port 515 nsew
rlabel metal1 s 5214 11430 5250 11771 4 vdd
port 515 nsew
rlabel metal1 s 222 19829 258 20170 4 vdd
port 515 nsew
rlabel metal1 s 7710 1160 7746 1501 4 vdd
port 515 nsew
rlabel metal1 s 4734 22989 4770 23330 4 vdd
port 515 nsew
rlabel metal1 s 18462 19829 18498 20170 4 vdd
port 515 nsew
rlabel metal1 s 5214 2449 5250 2790 4 vdd
port 515 nsew
rlabel metal1 s 16446 24569 16482 24910 4 vdd
port 515 nsew
rlabel metal1 s 10974 869 11010 1210 4 vdd
port 515 nsew
rlabel metal1 s 17214 24569 17250 24910 4 vdd
port 515 nsew
rlabel metal1 s 12702 15089 12738 15430 4 vdd
port 515 nsew
rlabel metal1 s 8958 18249 8994 18590 4 vdd
port 515 nsew
rlabel metal1 s 10206 16960 10242 17301 4 vdd
port 515 nsew
rlabel metal1 s 8478 7189 8514 7530 4 vdd
port 515 nsew
rlabel metal1 s 6462 16170 6498 16511 4 vdd
port 515 nsew
rlabel metal1 s 7230 13800 7266 14141 4 vdd
port 515 nsew
rlabel metal1 s 15966 18249 16002 18590 4 vdd
port 515 nsew
rlabel metal1 s 10206 23779 10242 24120 4 vdd
port 515 nsew
rlabel metal1 s 15966 5900 16002 6241 4 vdd
port 515 nsew
rlabel metal1 s 7230 19829 7266 20170 4 vdd
port 515 nsew
rlabel metal1 s 5982 10640 6018 10981 4 vdd
port 515 nsew
rlabel metal1 s 990 24569 1026 24910 4 vdd
port 515 nsew
rlabel metal1 s 10974 7979 11010 8320 4 vdd
port 515 nsew
rlabel metal1 s 3966 22199 4002 22540 4 vdd
port 515 nsew
rlabel metal1 s 12702 21700 12738 22041 4 vdd
port 515 nsew
rlabel metal1 s 8958 370 8994 711 4 vdd
port 515 nsew
rlabel metal1 s 4734 20619 4770 20960 4 vdd
port 515 nsew
rlabel metal1 s 15198 20619 15234 20960 4 vdd
port 515 nsew
rlabel metal1 s 10974 1160 11010 1501 4 vdd
port 515 nsew
rlabel metal1 s 2238 5110 2274 5451 4 vdd
port 515 nsew
rlabel metal1 s 8478 3530 8514 3871 4 vdd
port 515 nsew
rlabel metal1 s 13470 1160 13506 1501 4 vdd
port 515 nsew
rlabel metal1 s 2718 7189 2754 7530 4 vdd
port 515 nsew
rlabel metal1 s 5982 6690 6018 7031 4 vdd
port 515 nsew
rlabel metal1 s 12702 6399 12738 6740 4 vdd
port 515 nsew
rlabel metal1 s 222 16960 258 17301 4 vdd
port 515 nsew
rlabel metal1 s 12222 17459 12258 17800 4 vdd
port 515 nsew
rlabel metal1 s 7230 6399 7266 6740 4 vdd
port 515 nsew
rlabel metal1 s 3486 13010 3522 13351 4 vdd
port 515 nsew
rlabel metal1 s 19710 24860 19746 25201 4 vdd
port 515 nsew
rlabel metal1 s 3486 7189 3522 7530 4 vdd
port 515 nsew
rlabel metal1 s 13470 13010 13506 13351 4 vdd
port 515 nsew
rlabel metal1 s 8478 1659 8514 2000 4 vdd
port 515 nsew
rlabel metal1 s 5982 6399 6018 6740 4 vdd
port 515 nsew
rlabel metal1 s 1470 13800 1506 14141 4 vdd
port 515 nsew
rlabel metal1 s 13950 11430 13986 11771 4 vdd
port 515 nsew
rlabel metal1 s 1470 15380 1506 15721 4 vdd
port 515 nsew
rlabel metal1 s 8958 13800 8994 14141 4 vdd
port 515 nsew
rlabel metal1 s 7710 12719 7746 13060 4 vdd
port 515 nsew
rlabel metal1 s 7710 8270 7746 8611 4 vdd
port 515 nsew
rlabel metal1 s 8478 18540 8514 18881 4 vdd
port 515 nsew
rlabel metal1 s 10974 9060 11010 9401 4 vdd
port 515 nsew
rlabel metal1 s 12222 11929 12258 12270 4 vdd
port 515 nsew
rlabel metal1 s 5214 20910 5250 21251 4 vdd
port 515 nsew
rlabel metal1 s 14718 1659 14754 2000 4 vdd
port 515 nsew
rlabel metal1 s 12702 14299 12738 14640 4 vdd
port 515 nsew
rlabel metal1 s 15966 7979 16002 8320 4 vdd
port 515 nsew
rlabel metal1 s 222 13509 258 13850 4 vdd
port 515 nsew
rlabel metal1 s 10206 12719 10242 13060 4 vdd
port 515 nsew
rlabel metal1 s 14718 5900 14754 6241 4 vdd
port 515 nsew
rlabel metal1 s 4734 19039 4770 19380 4 vdd
port 515 nsew
rlabel metal1 s 19710 9850 19746 10191 4 vdd
port 515 nsew
rlabel metal1 s 8958 24860 8994 25201 4 vdd
port 515 nsew
rlabel metal1 s 1470 21700 1506 22041 4 vdd
port 515 nsew
rlabel metal1 s 13470 2740 13506 3081 4 vdd
port 515 nsew
rlabel metal1 s 5214 23779 5250 24120 4 vdd
port 515 nsew
rlabel metal1 s 15198 21409 15234 21750 4 vdd
port 515 nsew
rlabel metal1 s 4734 370 4770 711 4 vdd
port 515 nsew
rlabel metal1 s 18942 20120 18978 20461 4 vdd
port 515 nsew
rlabel metal1 s 7230 370 7266 711 4 vdd
port 515 nsew
rlabel metal1 s 10206 9060 10242 9401 4 vdd
port 515 nsew
rlabel metal1 s 18942 15879 18978 16220 4 vdd
port 515 nsew
rlabel metal1 s 15198 11139 15234 11480 4 vdd
port 515 nsew
rlabel metal1 s 1470 24860 1506 25201 4 vdd
port 515 nsew
rlabel metal1 s 7710 869 7746 1210 4 vdd
port 515 nsew
rlabel metal1 s 2238 3530 2274 3871 4 vdd
port 515 nsew
rlabel metal1 s 17694 24569 17730 24910 4 vdd
port 515 nsew
rlabel metal1 s 8958 12220 8994 12561 4 vdd
port 515 nsew
rlabel metal1 s 2238 1950 2274 2291 4 vdd
port 515 nsew
rlabel metal1 s 5214 16669 5250 17010 4 vdd
port 515 nsew
rlabel metal1 s 990 5900 1026 6241 4 vdd
port 515 nsew
rlabel metal1 s 3486 1950 3522 2291 4 vdd
port 515 nsew
rlabel metal1 s 10974 24569 11010 24910 4 vdd
port 515 nsew
rlabel metal1 s 3486 4029 3522 4370 4 vdd
port 515 nsew
rlabel metal1 s 14718 13010 14754 13351 4 vdd
port 515 nsew
rlabel metal1 s 222 20910 258 21251 4 vdd
port 515 nsew
rlabel metal1 s 3486 5609 3522 5950 4 vdd
port 515 nsew
rlabel metal1 s 12222 19039 12258 19380 4 vdd
port 515 nsew
rlabel metal1 s 3486 2740 3522 3081 4 vdd
port 515 nsew
rlabel metal1 s 2238 10640 2274 10981 4 vdd
port 515 nsew
rlabel metal1 s 17694 7979 17730 8320 4 vdd
port 515 nsew
rlabel metal1 s 13470 79 13506 420 4 vdd
port 515 nsew
rlabel metal1 s 12702 10640 12738 10981 4 vdd
port 515 nsew
rlabel metal1 s 5214 3239 5250 3580 4 vdd
port 515 nsew
rlabel metal1 s 6462 2740 6498 3081 4 vdd
port 515 nsew
rlabel metal1 s 10206 79 10242 420 4 vdd
port 515 nsew
rlabel metal1 s 7710 13010 7746 13351 4 vdd
port 515 nsew
rlabel metal1 s 7710 9559 7746 9900 4 vdd
port 515 nsew
rlabel metal1 s 17694 22490 17730 22831 4 vdd
port 515 nsew
rlabel metal1 s 990 12719 1026 13060 4 vdd
port 515 nsew
rlabel metal1 s 7230 10640 7266 10981 4 vdd
port 515 nsew
rlabel metal1 s 15198 3239 15234 3580 4 vdd
port 515 nsew
rlabel metal1 s 3486 11929 3522 12270 4 vdd
port 515 nsew
rlabel metal1 s 990 21409 1026 21750 4 vdd
port 515 nsew
rlabel metal1 s 13470 11929 13506 12270 4 vdd
port 515 nsew
rlabel metal1 s 18942 2449 18978 2790 4 vdd
port 515 nsew
rlabel metal1 s 1470 1659 1506 2000 4 vdd
port 515 nsew
rlabel metal1 s 1470 24569 1506 24910 4 vdd
port 515 nsew
rlabel metal1 s 6462 9060 6498 9401 4 vdd
port 515 nsew
rlabel metal1 s 13470 18540 13506 18881 4 vdd
port 515 nsew
rlabel metal1 s 15198 22490 15234 22831 4 vdd
port 515 nsew
rlabel metal1 s 5982 15380 6018 15721 4 vdd
port 515 nsew
rlabel metal1 s 14718 1160 14754 1501 4 vdd
port 515 nsew
rlabel metal1 s 12702 10349 12738 10690 4 vdd
port 515 nsew
rlabel metal1 s 13470 22490 13506 22831 4 vdd
port 515 nsew
rlabel metal1 s 2238 869 2274 1210 4 vdd
port 515 nsew
rlabel metal1 s 2718 79 2754 420 4 vdd
port 515 nsew
rlabel metal1 s 15198 1950 15234 2291 4 vdd
port 515 nsew
rlabel metal1 s 17214 14299 17250 14640 4 vdd
port 515 nsew
rlabel metal1 s 18462 8270 18498 8611 4 vdd
port 515 nsew
rlabel metal1 s 8478 22989 8514 23330 4 vdd
port 515 nsew
rlabel metal1 s 15966 15089 16002 15430 4 vdd
port 515 nsew
rlabel metal1 s 7230 1160 7266 1501 4 vdd
port 515 nsew
rlabel metal1 s 990 23280 1026 23621 4 vdd
port 515 nsew
rlabel metal1 s 15966 10640 16002 10981 4 vdd
port 515 nsew
rlabel metal1 s 3486 9559 3522 9900 4 vdd
port 515 nsew
rlabel metal1 s 3486 14590 3522 14931 4 vdd
port 515 nsew
rlabel metal1 s 222 14590 258 14931 4 vdd
port 515 nsew
rlabel metal1 s 11454 1950 11490 2291 4 vdd
port 515 nsew
rlabel metal1 s 2718 2740 2754 3081 4 vdd
port 515 nsew
rlabel metal1 s 11454 7189 11490 7530 4 vdd
port 515 nsew
rlabel metal1 s 18462 16960 18498 17301 4 vdd
port 515 nsew
rlabel metal1 s 16446 20619 16482 20960 4 vdd
port 515 nsew
rlabel metal1 s 17694 20120 17730 20461 4 vdd
port 515 nsew
rlabel metal1 s 7230 6690 7266 7031 4 vdd
port 515 nsew
rlabel metal1 s 9726 1950 9762 2291 4 vdd
port 515 nsew
rlabel metal1 s 2238 2449 2274 2790 4 vdd
port 515 nsew
rlabel metal1 s 15966 4029 16002 4370 4 vdd
port 515 nsew
rlabel metal1 s 7710 4320 7746 4661 4 vdd
port 515 nsew
rlabel metal1 s 10974 5110 11010 5451 4 vdd
port 515 nsew
rlabel metal1 s 15198 6690 15234 7031 4 vdd
port 515 nsew
rlabel metal1 s 17214 17459 17250 17800 4 vdd
port 515 nsew
rlabel metal1 s 12222 18540 12258 18881 4 vdd
port 515 nsew
rlabel metal1 s 17694 13509 17730 13850 4 vdd
port 515 nsew
rlabel metal1 s 18462 18540 18498 18881 4 vdd
port 515 nsew
rlabel metal1 s 3486 13509 3522 13850 4 vdd
port 515 nsew
rlabel metal1 s 14718 7979 14754 8320 4 vdd
port 515 nsew
rlabel metal1 s 2718 22989 2754 23330 4 vdd
port 515 nsew
rlabel metal1 s 17694 21700 17730 22041 4 vdd
port 515 nsew
rlabel metal1 s 18942 16960 18978 17301 4 vdd
port 515 nsew
rlabel metal1 s 3966 11430 4002 11771 4 vdd
port 515 nsew
rlabel metal1 s 5982 4320 6018 4661 4 vdd
port 515 nsew
rlabel metal1 s 14718 23280 14754 23621 4 vdd
port 515 nsew
rlabel metal1 s 19710 5900 19746 6241 4 vdd
port 515 nsew
rlabel metal1 s 7230 21409 7266 21750 4 vdd
port 515 nsew
rlabel metal1 s 15198 19330 15234 19671 4 vdd
port 515 nsew
rlabel metal1 s 16446 13800 16482 14141 4 vdd
port 515 nsew
rlabel metal1 s 3486 22989 3522 23330 4 vdd
port 515 nsew
rlabel metal1 s 222 15380 258 15721 4 vdd
port 515 nsew
rlabel metal1 s 6462 13010 6498 13351 4 vdd
port 515 nsew
rlabel metal1 s 8478 8769 8514 9110 4 vdd
port 515 nsew
rlabel metal1 s 7710 16669 7746 17010 4 vdd
port 515 nsew
rlabel metal1 s 4734 7979 4770 8320 4 vdd
port 515 nsew
rlabel metal1 s 18462 18249 18498 18590 4 vdd
port 515 nsew
rlabel metal1 s 13470 19330 13506 19671 4 vdd
port 515 nsew
rlabel metal1 s 17694 17459 17730 17800 4 vdd
port 515 nsew
rlabel metal1 s 7230 16669 7266 17010 4 vdd
port 515 nsew
rlabel metal1 s 4734 10640 4770 10981 4 vdd
port 515 nsew
rlabel metal1 s 3966 1950 4002 2291 4 vdd
port 515 nsew
rlabel metal1 s 7710 7189 7746 7530 4 vdd
port 515 nsew
rlabel metal1 s 990 10640 1026 10981 4 vdd
port 515 nsew
rlabel metal1 s 9726 11430 9762 11771 4 vdd
port 515 nsew
rlabel metal1 s 7710 15089 7746 15430 4 vdd
port 515 nsew
rlabel metal1 s 2238 22989 2274 23330 4 vdd
port 515 nsew
rlabel metal1 s 8958 7480 8994 7821 4 vdd
port 515 nsew
rlabel metal1 s 9726 4819 9762 5160 4 vdd
port 515 nsew
rlabel metal1 s 6462 12220 6498 12561 4 vdd
port 515 nsew
rlabel metal1 s 18942 9559 18978 9900 4 vdd
port 515 nsew
rlabel metal1 s 9726 17459 9762 17800 4 vdd
port 515 nsew
rlabel metal1 s 17694 19330 17730 19671 4 vdd
port 515 nsew
rlabel metal1 s 7230 20619 7266 20960 4 vdd
port 515 nsew
rlabel metal1 s 14718 370 14754 711 4 vdd
port 515 nsew
rlabel metal1 s 3966 22490 4002 22831 4 vdd
port 515 nsew
rlabel metal1 s 2238 7480 2274 7821 4 vdd
port 515 nsew
rlabel metal1 s 4734 5110 4770 5451 4 vdd
port 515 nsew
rlabel metal1 s 6462 13800 6498 14141 4 vdd
port 515 nsew
rlabel metal1 s 8958 13509 8994 13850 4 vdd
port 515 nsew
rlabel metal1 s 1470 16669 1506 17010 4 vdd
port 515 nsew
rlabel metal1 s 14718 17459 14754 17800 4 vdd
port 515 nsew
rlabel metal1 s 5982 3239 6018 3580 4 vdd
port 515 nsew
rlabel metal1 s 16446 11139 16482 11480 4 vdd
port 515 nsew
rlabel metal1 s 990 2740 1026 3081 4 vdd
port 515 nsew
rlabel metal1 s 4734 13010 4770 13351 4 vdd
port 515 nsew
rlabel metal1 s 12222 5900 12258 6241 4 vdd
port 515 nsew
rlabel metal1 s 10974 7480 11010 7821 4 vdd
port 515 nsew
rlabel metal1 s 12702 19330 12738 19671 4 vdd
port 515 nsew
rlabel metal1 s 2238 19330 2274 19671 4 vdd
port 515 nsew
rlabel metal1 s 2238 8769 2274 9110 4 vdd
port 515 nsew
rlabel metal1 s 13950 1950 13986 2291 4 vdd
port 515 nsew
rlabel metal1 s 8958 20910 8994 21251 4 vdd
port 515 nsew
rlabel metal1 s 13950 869 13986 1210 4 vdd
port 515 nsew
rlabel metal1 s 19710 7979 19746 8320 4 vdd
port 515 nsew
rlabel metal1 s 10974 14299 11010 14640 4 vdd
port 515 nsew
rlabel metal1 s 2718 18249 2754 18590 4 vdd
port 515 nsew
rlabel metal1 s 2718 7480 2754 7821 4 vdd
port 515 nsew
rlabel metal1 s 8958 2449 8994 2790 4 vdd
port 515 nsew
rlabel metal1 s 8958 22490 8994 22831 4 vdd
port 515 nsew
rlabel metal1 s 10974 15089 11010 15430 4 vdd
port 515 nsew
rlabel metal1 s 14718 9060 14754 9401 4 vdd
port 515 nsew
rlabel metal1 s 11454 5110 11490 5451 4 vdd
port 515 nsew
rlabel metal1 s 12222 5110 12258 5451 4 vdd
port 515 nsew
rlabel metal1 s 14718 9559 14754 9900 4 vdd
port 515 nsew
rlabel metal1 s 3966 23280 4002 23621 4 vdd
port 515 nsew
rlabel metal1 s 14718 2740 14754 3081 4 vdd
port 515 nsew
rlabel metal1 s 15198 18540 15234 18881 4 vdd
port 515 nsew
rlabel metal1 s 3966 5900 4002 6241 4 vdd
port 515 nsew
rlabel metal1 s 7710 17459 7746 17800 4 vdd
port 515 nsew
rlabel metal1 s 12702 13509 12738 13850 4 vdd
port 515 nsew
rlabel metal1 s 17214 2449 17250 2790 4 vdd
port 515 nsew
rlabel metal1 s 18462 17459 18498 17800 4 vdd
port 515 nsew
rlabel metal1 s 222 23280 258 23621 4 vdd
port 515 nsew
rlabel metal1 s 12702 16669 12738 17010 4 vdd
port 515 nsew
rlabel metal1 s 15966 21409 16002 21750 4 vdd
port 515 nsew
rlabel metal1 s 16446 7480 16482 7821 4 vdd
port 515 nsew
rlabel metal1 s 13950 22490 13986 22831 4 vdd
port 515 nsew
rlabel metal1 s 13950 370 13986 711 4 vdd
port 515 nsew
rlabel metal1 s 8478 9559 8514 9900 4 vdd
port 515 nsew
rlabel metal1 s 7710 14299 7746 14640 4 vdd
port 515 nsew
rlabel metal1 s 9726 9060 9762 9401 4 vdd
port 515 nsew
rlabel metal1 s 8478 5900 8514 6241 4 vdd
port 515 nsew
rlabel metal1 s 8958 12719 8994 13060 4 vdd
port 515 nsew
rlabel metal1 s 222 8769 258 9110 4 vdd
port 515 nsew
rlabel metal1 s 222 14299 258 14640 4 vdd
port 515 nsew
rlabel metal1 s 990 22490 1026 22831 4 vdd
port 515 nsew
rlabel metal1 s 8478 11929 8514 12270 4 vdd
port 515 nsew
rlabel metal1 s 13470 17750 13506 18091 4 vdd
port 515 nsew
rlabel metal1 s 18942 1659 18978 2000 4 vdd
port 515 nsew
rlabel metal1 s 17694 3239 17730 3580 4 vdd
port 515 nsew
rlabel metal1 s 222 3530 258 3871 4 vdd
port 515 nsew
rlabel metal1 s 3966 7979 4002 8320 4 vdd
port 515 nsew
rlabel metal1 s 18942 19829 18978 20170 4 vdd
port 515 nsew
rlabel metal1 s 11454 13509 11490 13850 4 vdd
port 515 nsew
rlabel metal1 s 8478 8270 8514 8611 4 vdd
port 515 nsew
rlabel metal1 s 4734 19330 4770 19671 4 vdd
port 515 nsew
rlabel metal1 s 8478 2449 8514 2790 4 vdd
port 515 nsew
rlabel metal1 s 19710 12719 19746 13060 4 vdd
port 515 nsew
rlabel metal1 s 6462 8769 6498 9110 4 vdd
port 515 nsew
rlabel metal1 s 9726 4320 9762 4661 4 vdd
port 515 nsew
rlabel metal1 s 10974 1950 11010 2291 4 vdd
port 515 nsew
rlabel metal1 s 222 11139 258 11480 4 vdd
port 515 nsew
rlabel metal1 s 1470 7189 1506 7530 4 vdd
port 515 nsew
rlabel metal1 s 13470 4320 13506 4661 4 vdd
port 515 nsew
rlabel metal1 s 16446 17459 16482 17800 4 vdd
port 515 nsew
rlabel metal1 s 15198 6399 15234 6740 4 vdd
port 515 nsew
rlabel metal1 s 5982 24070 6018 24411 4 vdd
port 515 nsew
rlabel metal1 s 18462 21700 18498 22041 4 vdd
port 515 nsew
rlabel metal1 s 6462 13509 6498 13850 4 vdd
port 515 nsew
rlabel metal1 s 18942 8769 18978 9110 4 vdd
port 515 nsew
rlabel metal1 s 19710 15879 19746 16220 4 vdd
port 515 nsew
rlabel metal1 s 11454 9850 11490 10191 4 vdd
port 515 nsew
rlabel metal1 s 16446 24070 16482 24411 4 vdd
port 515 nsew
rlabel metal1 s 990 21700 1026 22041 4 vdd
port 515 nsew
rlabel metal1 s 3486 12220 3522 12561 4 vdd
port 515 nsew
rlabel metal1 s 12222 1659 12258 2000 4 vdd
port 515 nsew
rlabel metal1 s 8958 22989 8994 23330 4 vdd
port 515 nsew
rlabel metal1 s 17214 2740 17250 3081 4 vdd
port 515 nsew
rlabel metal1 s 18942 9060 18978 9401 4 vdd
port 515 nsew
rlabel metal1 s 6462 7480 6498 7821 4 vdd
port 515 nsew
rlabel metal1 s 18462 1950 18498 2291 4 vdd
port 515 nsew
rlabel metal1 s 12222 4029 12258 4370 4 vdd
port 515 nsew
rlabel metal1 s 17214 8769 17250 9110 4 vdd
port 515 nsew
rlabel metal1 s 3966 4029 4002 4370 4 vdd
port 515 nsew
rlabel metal1 s 17694 24860 17730 25201 4 vdd
port 515 nsew
rlabel metal1 s 1470 3530 1506 3871 4 vdd
port 515 nsew
rlabel metal1 s 5982 7189 6018 7530 4 vdd
port 515 nsew
rlabel metal1 s 11454 10349 11490 10690 4 vdd
port 515 nsew
rlabel metal1 s 10206 13010 10242 13351 4 vdd
port 515 nsew
rlabel metal1 s 222 18249 258 18590 4 vdd
port 515 nsew
rlabel metal1 s 1470 11929 1506 12270 4 vdd
port 515 nsew
rlabel metal1 s 10206 20120 10242 20461 4 vdd
port 515 nsew
rlabel metal1 s 5982 2740 6018 3081 4 vdd
port 515 nsew
rlabel metal1 s 13470 13509 13506 13850 4 vdd
port 515 nsew
rlabel metal1 s 16446 15879 16482 16220 4 vdd
port 515 nsew
rlabel metal1 s 2718 7979 2754 8320 4 vdd
port 515 nsew
rlabel metal1 s 18942 23280 18978 23621 4 vdd
port 515 nsew
rlabel metal1 s 990 370 1026 711 4 vdd
port 515 nsew
rlabel metal1 s 5214 24569 5250 24910 4 vdd
port 515 nsew
rlabel metal1 s 8958 20619 8994 20960 4 vdd
port 515 nsew
rlabel metal1 s 18462 869 18498 1210 4 vdd
port 515 nsew
rlabel metal1 s 2238 22490 2274 22831 4 vdd
port 515 nsew
rlabel metal1 s 9726 16170 9762 16511 4 vdd
port 515 nsew
rlabel metal1 s 3966 12220 4002 12561 4 vdd
port 515 nsew
rlabel metal1 s 8478 79 8514 420 4 vdd
port 515 nsew
rlabel metal1 s 18942 4320 18978 4661 4 vdd
port 515 nsew
rlabel metal1 s 3486 15380 3522 15721 4 vdd
port 515 nsew
rlabel metal1 s 12222 9060 12258 9401 4 vdd
port 515 nsew
rlabel metal1 s 16446 7979 16482 8320 4 vdd
port 515 nsew
rlabel metal1 s 9726 19330 9762 19671 4 vdd
port 515 nsew
rlabel metal1 s 6462 5900 6498 6241 4 vdd
port 515 nsew
rlabel metal1 s 18462 21409 18498 21750 4 vdd
port 515 nsew
rlabel metal1 s 8958 15089 8994 15430 4 vdd
port 515 nsew
rlabel metal1 s 2238 20619 2274 20960 4 vdd
port 515 nsew
rlabel metal1 s 6462 20120 6498 20461 4 vdd
port 515 nsew
rlabel metal1 s 12702 3530 12738 3871 4 vdd
port 515 nsew
rlabel metal1 s 18942 21409 18978 21750 4 vdd
port 515 nsew
rlabel metal1 s 17214 10349 17250 10690 4 vdd
port 515 nsew
rlabel metal1 s 17694 13800 17730 14141 4 vdd
port 515 nsew
rlabel metal1 s 13950 18540 13986 18881 4 vdd
port 515 nsew
rlabel metal1 s 990 13010 1026 13351 4 vdd
port 515 nsew
rlabel metal1 s 17214 869 17250 1210 4 vdd
port 515 nsew
rlabel metal1 s 10974 15879 11010 16220 4 vdd
port 515 nsew
rlabel metal1 s 11454 3239 11490 3580 4 vdd
port 515 nsew
rlabel metal1 s 12702 24070 12738 24411 4 vdd
port 515 nsew
rlabel metal1 s 18942 10349 18978 10690 4 vdd
port 515 nsew
rlabel metal1 s 15198 23779 15234 24120 4 vdd
port 515 nsew
rlabel metal1 s 18942 11929 18978 12270 4 vdd
port 515 nsew
rlabel metal1 s 3486 5110 3522 5451 4 vdd
port 515 nsew
rlabel metal1 s 17214 12719 17250 13060 4 vdd
port 515 nsew
rlabel metal1 s 15966 20910 16002 21251 4 vdd
port 515 nsew
rlabel metal1 s 16446 18540 16482 18881 4 vdd
port 515 nsew
rlabel metal1 s 4734 2740 4770 3081 4 vdd
port 515 nsew
rlabel metal1 s 17694 16669 17730 17010 4 vdd
port 515 nsew
rlabel metal1 s 8958 23280 8994 23621 4 vdd
port 515 nsew
rlabel metal1 s 4734 23280 4770 23621 4 vdd
port 515 nsew
rlabel metal1 s 1470 11139 1506 11480 4 vdd
port 515 nsew
rlabel metal1 s 17694 10349 17730 10690 4 vdd
port 515 nsew
rlabel metal1 s 12222 8769 12258 9110 4 vdd
port 515 nsew
rlabel metal1 s 14718 4029 14754 4370 4 vdd
port 515 nsew
rlabel metal1 s 14718 4819 14754 5160 4 vdd
port 515 nsew
rlabel metal1 s 10206 7979 10242 8320 4 vdd
port 515 nsew
rlabel metal1 s 10974 21409 11010 21750 4 vdd
port 515 nsew
rlabel metal1 s 14718 19330 14754 19671 4 vdd
port 515 nsew
rlabel metal1 s 17214 14590 17250 14931 4 vdd
port 515 nsew
rlabel metal1 s 16446 21409 16482 21750 4 vdd
port 515 nsew
rlabel metal1 s 8478 19829 8514 20170 4 vdd
port 515 nsew
rlabel metal1 s 5982 14299 6018 14640 4 vdd
port 515 nsew
rlabel metal1 s 15198 11430 15234 11771 4 vdd
port 515 nsew
rlabel metal1 s 15966 5609 16002 5950 4 vdd
port 515 nsew
rlabel metal1 s 13950 8270 13986 8611 4 vdd
port 515 nsew
rlabel metal1 s 2238 11430 2274 11771 4 vdd
port 515 nsew
rlabel metal1 s 10974 9559 11010 9900 4 vdd
port 515 nsew
rlabel metal1 s 18462 15879 18498 16220 4 vdd
port 515 nsew
rlabel metal1 s 7710 13509 7746 13850 4 vdd
port 515 nsew
rlabel metal1 s 12222 12719 12258 13060 4 vdd
port 515 nsew
rlabel metal1 s 11454 15879 11490 16220 4 vdd
port 515 nsew
rlabel metal1 s 12702 11430 12738 11771 4 vdd
port 515 nsew
rlabel metal1 s 3486 8769 3522 9110 4 vdd
port 515 nsew
rlabel metal1 s 8958 5110 8994 5451 4 vdd
port 515 nsew
rlabel metal1 s 990 4320 1026 4661 4 vdd
port 515 nsew
rlabel metal1 s 13470 21700 13506 22041 4 vdd
port 515 nsew
rlabel metal1 s 13950 3530 13986 3871 4 vdd
port 515 nsew
rlabel metal1 s 14718 19829 14754 20170 4 vdd
port 515 nsew
rlabel metal1 s 15966 7189 16002 7530 4 vdd
port 515 nsew
rlabel metal1 s 7710 79 7746 420 4 vdd
port 515 nsew
rlabel metal1 s 7710 6690 7746 7031 4 vdd
port 515 nsew
rlabel metal1 s 10974 22490 11010 22831 4 vdd
port 515 nsew
rlabel metal1 s 7710 19039 7746 19380 4 vdd
port 515 nsew
rlabel metal1 s 4734 24860 4770 25201 4 vdd
port 515 nsew
rlabel metal1 s 19710 14299 19746 14640 4 vdd
port 515 nsew
rlabel metal1 s 13950 11139 13986 11480 4 vdd
port 515 nsew
rlabel metal1 s 6462 15879 6498 16220 4 vdd
port 515 nsew
rlabel metal1 s 13470 8270 13506 8611 4 vdd
port 515 nsew
rlabel metal1 s 1470 2449 1506 2790 4 vdd
port 515 nsew
rlabel metal1 s 990 11929 1026 12270 4 vdd
port 515 nsew
rlabel metal1 s 15198 4029 15234 4370 4 vdd
port 515 nsew
rlabel metal1 s 18462 370 18498 711 4 vdd
port 515 nsew
rlabel metal1 s 5214 7979 5250 8320 4 vdd
port 515 nsew
rlabel metal1 s 7230 7979 7266 8320 4 vdd
port 515 nsew
rlabel metal1 s 15198 19039 15234 19380 4 vdd
port 515 nsew
rlabel metal1 s 7710 18540 7746 18881 4 vdd
port 515 nsew
rlabel metal1 s 15198 11929 15234 12270 4 vdd
port 515 nsew
rlabel metal1 s 16446 23779 16482 24120 4 vdd
port 515 nsew
rlabel metal1 s 4734 15380 4770 15721 4 vdd
port 515 nsew
rlabel metal1 s 7710 3239 7746 3580 4 vdd
port 515 nsew
rlabel metal1 s 18942 17750 18978 18091 4 vdd
port 515 nsew
rlabel metal1 s 11454 4029 11490 4370 4 vdd
port 515 nsew
rlabel metal1 s 6462 24569 6498 24910 4 vdd
port 515 nsew
rlabel metal1 s 222 9559 258 9900 4 vdd
port 515 nsew
rlabel metal1 s 10206 13509 10242 13850 4 vdd
port 515 nsew
rlabel metal1 s 14718 5609 14754 5950 4 vdd
port 515 nsew
rlabel metal1 s 8958 17459 8994 17800 4 vdd
port 515 nsew
rlabel metal1 s 19710 1160 19746 1501 4 vdd
port 515 nsew
rlabel metal1 s 12702 5609 12738 5950 4 vdd
port 515 nsew
rlabel metal1 s 2238 10349 2274 10690 4 vdd
port 515 nsew
rlabel metal1 s 17214 18249 17250 18590 4 vdd
port 515 nsew
rlabel metal1 s 18462 23280 18498 23621 4 vdd
port 515 nsew
rlabel metal1 s 3486 22490 3522 22831 4 vdd
port 515 nsew
rlabel metal1 s 9726 1659 9762 2000 4 vdd
port 515 nsew
rlabel metal1 s 10206 3530 10242 3871 4 vdd
port 515 nsew
rlabel metal1 s 990 15380 1026 15721 4 vdd
port 515 nsew
rlabel metal1 s 12222 79 12258 420 4 vdd
port 515 nsew
rlabel metal1 s 8478 20619 8514 20960 4 vdd
port 515 nsew
rlabel metal1 s 13470 8769 13506 9110 4 vdd
port 515 nsew
rlabel metal1 s 5982 13509 6018 13850 4 vdd
port 515 nsew
rlabel metal1 s 14718 10349 14754 10690 4 vdd
port 515 nsew
rlabel metal1 s 5982 13800 6018 14141 4 vdd
port 515 nsew
rlabel metal1 s 3486 18249 3522 18590 4 vdd
port 515 nsew
rlabel metal1 s 17214 1950 17250 2291 4 vdd
port 515 nsew
rlabel metal1 s 19710 13509 19746 13850 4 vdd
port 515 nsew
rlabel metal1 s 5214 6399 5250 6740 4 vdd
port 515 nsew
rlabel metal1 s 10974 2740 11010 3081 4 vdd
port 515 nsew
rlabel metal1 s 5214 24860 5250 25201 4 vdd
port 515 nsew
rlabel metal1 s 9726 9850 9762 10191 4 vdd
port 515 nsew
rlabel metal1 s 16446 13010 16482 13351 4 vdd
port 515 nsew
rlabel metal1 s 2718 5609 2754 5950 4 vdd
port 515 nsew
rlabel metal1 s 3486 16669 3522 17010 4 vdd
port 515 nsew
rlabel metal1 s 7230 16960 7266 17301 4 vdd
port 515 nsew
rlabel metal1 s 11454 19829 11490 20170 4 vdd
port 515 nsew
rlabel metal1 s 15966 22490 16002 22831 4 vdd
port 515 nsew
rlabel metal1 s 12222 4320 12258 4661 4 vdd
port 515 nsew
rlabel metal1 s 3486 20120 3522 20461 4 vdd
port 515 nsew
rlabel metal1 s 9726 24569 9762 24910 4 vdd
port 515 nsew
rlabel metal1 s 1470 4029 1506 4370 4 vdd
port 515 nsew
rlabel metal1 s 17694 370 17730 711 4 vdd
port 515 nsew
rlabel metal1 s 19710 18249 19746 18590 4 vdd
port 515 nsew
rlabel metal1 s 990 1659 1026 2000 4 vdd
port 515 nsew
rlabel metal1 s 12222 16669 12258 17010 4 vdd
port 515 nsew
rlabel metal1 s 2238 14590 2274 14931 4 vdd
port 515 nsew
rlabel metal1 s 12702 20120 12738 20461 4 vdd
port 515 nsew
rlabel metal1 s 6462 16669 6498 17010 4 vdd
port 515 nsew
rlabel metal1 s 6462 1950 6498 2291 4 vdd
port 515 nsew
rlabel metal1 s 11454 2740 11490 3081 4 vdd
port 515 nsew
rlabel metal1 s 12702 9559 12738 9900 4 vdd
port 515 nsew
rlabel metal1 s 17214 19330 17250 19671 4 vdd
port 515 nsew
rlabel metal1 s 2238 9850 2274 10191 4 vdd
port 515 nsew
rlabel metal1 s 9726 11139 9762 11480 4 vdd
port 515 nsew
rlabel metal1 s 4734 11430 4770 11771 4 vdd
port 515 nsew
rlabel metal1 s 13470 15879 13506 16220 4 vdd
port 515 nsew
rlabel metal1 s 8958 16669 8994 17010 4 vdd
port 515 nsew
rlabel metal1 s 14718 6690 14754 7031 4 vdd
port 515 nsew
rlabel metal1 s 7710 11139 7746 11480 4 vdd
port 515 nsew
rlabel metal1 s 10974 24860 11010 25201 4 vdd
port 515 nsew
rlabel metal1 s 4734 7480 4770 7821 4 vdd
port 515 nsew
rlabel metal1 s 15198 2449 15234 2790 4 vdd
port 515 nsew
rlabel metal1 s 7710 4029 7746 4370 4 vdd
port 515 nsew
rlabel metal1 s 8478 19039 8514 19380 4 vdd
port 515 nsew
rlabel metal1 s 1470 10640 1506 10981 4 vdd
port 515 nsew
rlabel metal1 s 2718 23779 2754 24120 4 vdd
port 515 nsew
rlabel metal1 s 8478 12719 8514 13060 4 vdd
port 515 nsew
rlabel metal1 s 18942 14590 18978 14931 4 vdd
port 515 nsew
rlabel metal1 s 3966 3239 4002 3580 4 vdd
port 515 nsew
rlabel metal1 s 4734 18540 4770 18881 4 vdd
port 515 nsew
rlabel metal1 s 8478 2740 8514 3081 4 vdd
port 515 nsew
rlabel metal1 s 11454 17750 11490 18091 4 vdd
port 515 nsew
rlabel metal1 s 2238 21700 2274 22041 4 vdd
port 515 nsew
rlabel metal1 s 19710 9559 19746 9900 4 vdd
port 515 nsew
rlabel metal1 s 7710 370 7746 711 4 vdd
port 515 nsew
rlabel metal1 s 8958 14299 8994 14640 4 vdd
port 515 nsew
rlabel metal1 s 5982 15879 6018 16220 4 vdd
port 515 nsew
rlabel metal1 s 15198 9559 15234 9900 4 vdd
port 515 nsew
rlabel metal1 s 5214 13010 5250 13351 4 vdd
port 515 nsew
rlabel metal1 s 11454 9559 11490 9900 4 vdd
port 515 nsew
rlabel metal1 s 13950 14590 13986 14931 4 vdd
port 515 nsew
rlabel metal1 s 9726 8270 9762 8611 4 vdd
port 515 nsew
rlabel metal1 s 13950 6690 13986 7031 4 vdd
port 515 nsew
rlabel metal1 s 5982 4819 6018 5160 4 vdd
port 515 nsew
rlabel metal1 s 13950 23779 13986 24120 4 vdd
port 515 nsew
rlabel metal1 s 5214 12220 5250 12561 4 vdd
port 515 nsew
rlabel metal1 s 7230 16170 7266 16511 4 vdd
port 515 nsew
rlabel metal1 s 9726 6399 9762 6740 4 vdd
port 515 nsew
rlabel metal1 s 990 1950 1026 2291 4 vdd
port 515 nsew
rlabel metal1 s 9726 5609 9762 5950 4 vdd
port 515 nsew
rlabel metal1 s 6462 24070 6498 24411 4 vdd
port 515 nsew
rlabel metal1 s 2718 15380 2754 15721 4 vdd
port 515 nsew
rlabel metal1 s 12222 19330 12258 19671 4 vdd
port 515 nsew
rlabel metal1 s 17214 9850 17250 10191 4 vdd
port 515 nsew
rlabel metal1 s 2718 12220 2754 12561 4 vdd
port 515 nsew
rlabel metal1 s 4734 6399 4770 6740 4 vdd
port 515 nsew
rlabel metal1 s 17214 6690 17250 7031 4 vdd
port 515 nsew
rlabel metal1 s 222 23779 258 24120 4 vdd
port 515 nsew
rlabel metal1 s 17694 17750 17730 18091 4 vdd
port 515 nsew
rlabel metal1 s 14718 4320 14754 4661 4 vdd
port 515 nsew
rlabel metal1 s 5214 23280 5250 23621 4 vdd
port 515 nsew
rlabel metal1 s 1470 15879 1506 16220 4 vdd
port 515 nsew
rlabel metal1 s 5982 24860 6018 25201 4 vdd
port 515 nsew
rlabel metal1 s 5214 4819 5250 5160 4 vdd
port 515 nsew
rlabel metal1 s 10206 5609 10242 5950 4 vdd
port 515 nsew
rlabel metal1 s 18942 9850 18978 10191 4 vdd
port 515 nsew
rlabel metal1 s 3486 7480 3522 7821 4 vdd
port 515 nsew
rlabel metal1 s 222 21409 258 21750 4 vdd
port 515 nsew
rlabel metal1 s 3966 6690 4002 7031 4 vdd
port 515 nsew
rlabel metal1 s 6462 17750 6498 18091 4 vdd
port 515 nsew
rlabel metal1 s 18942 21700 18978 22041 4 vdd
port 515 nsew
rlabel metal1 s 5982 10349 6018 10690 4 vdd
port 515 nsew
rlabel metal1 s 15198 5900 15234 6241 4 vdd
port 515 nsew
rlabel metal1 s 10206 17459 10242 17800 4 vdd
port 515 nsew
rlabel metal1 s 6462 21700 6498 22041 4 vdd
port 515 nsew
rlabel metal1 s 3486 19039 3522 19380 4 vdd
port 515 nsew
rlabel metal1 s 15966 869 16002 1210 4 vdd
port 515 nsew
rlabel metal1 s 19710 8769 19746 9110 4 vdd
port 515 nsew
rlabel metal1 s 18462 12220 18498 12561 4 vdd
port 515 nsew
rlabel metal1 s 1470 8769 1506 9110 4 vdd
port 515 nsew
rlabel metal1 s 7710 21409 7746 21750 4 vdd
port 515 nsew
rlabel metal1 s 2718 17459 2754 17800 4 vdd
port 515 nsew
rlabel metal1 s 12222 7480 12258 7821 4 vdd
port 515 nsew
rlabel metal1 s 2238 4819 2274 5160 4 vdd
port 515 nsew
rlabel metal1 s 11454 2449 11490 2790 4 vdd
port 515 nsew
rlabel metal1 s 1470 6399 1506 6740 4 vdd
port 515 nsew
rlabel metal1 s 5214 5900 5250 6241 4 vdd
port 515 nsew
rlabel metal1 s 13950 13800 13986 14141 4 vdd
port 515 nsew
rlabel metal1 s 17214 9559 17250 9900 4 vdd
port 515 nsew
rlabel metal1 s 8958 22199 8994 22540 4 vdd
port 515 nsew
rlabel metal1 s 15198 23280 15234 23621 4 vdd
port 515 nsew
rlabel metal1 s 16446 11430 16482 11771 4 vdd
port 515 nsew
rlabel metal1 s 17214 18540 17250 18881 4 vdd
port 515 nsew
rlabel metal1 s 17214 17750 17250 18091 4 vdd
port 515 nsew
rlabel metal1 s 12702 7979 12738 8320 4 vdd
port 515 nsew
rlabel metal1 s 13950 9060 13986 9401 4 vdd
port 515 nsew
rlabel metal1 s 7230 7189 7266 7530 4 vdd
port 515 nsew
rlabel metal1 s 12702 2740 12738 3081 4 vdd
port 515 nsew
rlabel metal1 s 14718 11929 14754 12270 4 vdd
port 515 nsew
rlabel metal1 s 10206 16170 10242 16511 4 vdd
port 515 nsew
rlabel metal1 s 10206 10640 10242 10981 4 vdd
port 515 nsew
rlabel metal1 s 3486 4819 3522 5160 4 vdd
port 515 nsew
rlabel metal1 s 18942 22199 18978 22540 4 vdd
port 515 nsew
rlabel metal1 s 19710 7189 19746 7530 4 vdd
port 515 nsew
rlabel metal1 s 7710 17750 7746 18091 4 vdd
port 515 nsew
rlabel metal1 s 13470 16669 13506 17010 4 vdd
port 515 nsew
rlabel metal1 s 7230 2740 7266 3081 4 vdd
port 515 nsew
rlabel metal1 s 2718 13010 2754 13351 4 vdd
port 515 nsew
rlabel metal1 s 18942 11430 18978 11771 4 vdd
port 515 nsew
rlabel metal1 s 10206 11929 10242 12270 4 vdd
port 515 nsew
rlabel metal1 s 7230 3239 7266 3580 4 vdd
port 515 nsew
rlabel metal1 s 11454 16170 11490 16511 4 vdd
port 515 nsew
rlabel metal1 s 13470 1950 13506 2291 4 vdd
port 515 nsew
rlabel metal1 s 17694 2449 17730 2790 4 vdd
port 515 nsew
rlabel metal1 s 13950 6399 13986 6740 4 vdd
port 515 nsew
rlabel metal1 s 3966 16669 4002 17010 4 vdd
port 515 nsew
rlabel metal1 s 13470 20619 13506 20960 4 vdd
port 515 nsew
rlabel metal1 s 17214 24860 17250 25201 4 vdd
port 515 nsew
rlabel metal1 s 2718 6399 2754 6740 4 vdd
port 515 nsew
rlabel metal1 s 10206 17750 10242 18091 4 vdd
port 515 nsew
rlabel metal1 s 16446 17750 16482 18091 4 vdd
port 515 nsew
rlabel metal1 s 2718 1659 2754 2000 4 vdd
port 515 nsew
rlabel metal1 s 19710 1950 19746 2291 4 vdd
port 515 nsew
rlabel metal1 s 19710 11430 19746 11771 4 vdd
port 515 nsew
rlabel metal1 s 7710 7979 7746 8320 4 vdd
port 515 nsew
rlabel metal1 s 14718 21700 14754 22041 4 vdd
port 515 nsew
rlabel metal1 s 8958 11430 8994 11771 4 vdd
port 515 nsew
rlabel metal1 s 2718 11430 2754 11771 4 vdd
port 515 nsew
rlabel metal1 s 12702 16960 12738 17301 4 vdd
port 515 nsew
rlabel metal1 s 10206 20910 10242 21251 4 vdd
port 515 nsew
rlabel metal1 s 990 9559 1026 9900 4 vdd
port 515 nsew
rlabel metal1 s 10206 20619 10242 20960 4 vdd
port 515 nsew
rlabel metal1 s 4734 20120 4770 20461 4 vdd
port 515 nsew
rlabel metal1 s 1470 3239 1506 3580 4 vdd
port 515 nsew
rlabel metal1 s 8958 9060 8994 9401 4 vdd
port 515 nsew
rlabel metal1 s 9726 7979 9762 8320 4 vdd
port 515 nsew
rlabel metal1 s 8478 11139 8514 11480 4 vdd
port 515 nsew
rlabel metal1 s 7710 22989 7746 23330 4 vdd
port 515 nsew
rlabel metal1 s 6462 15089 6498 15430 4 vdd
port 515 nsew
rlabel metal1 s 222 16669 258 17010 4 vdd
port 515 nsew
rlabel metal1 s 5982 8270 6018 8611 4 vdd
port 515 nsew
rlabel metal1 s 7230 3530 7266 3871 4 vdd
port 515 nsew
rlabel metal1 s 8958 16960 8994 17301 4 vdd
port 515 nsew
rlabel metal1 s 16446 6399 16482 6740 4 vdd
port 515 nsew
rlabel metal1 s 15966 11929 16002 12270 4 vdd
port 515 nsew
rlabel metal1 s 990 16170 1026 16511 4 vdd
port 515 nsew
rlabel metal1 s 7230 14590 7266 14931 4 vdd
port 515 nsew
rlabel metal1 s 5214 13509 5250 13850 4 vdd
port 515 nsew
rlabel metal1 s 2718 20619 2754 20960 4 vdd
port 515 nsew
rlabel metal1 s 5214 24070 5250 24411 4 vdd
port 515 nsew
rlabel metal1 s 12222 9850 12258 10191 4 vdd
port 515 nsew
rlabel metal1 s 13950 16960 13986 17301 4 vdd
port 515 nsew
rlabel metal1 s 10974 23280 11010 23621 4 vdd
port 515 nsew
rlabel metal1 s 14718 16170 14754 16511 4 vdd
port 515 nsew
rlabel metal1 s 19710 15089 19746 15430 4 vdd
port 515 nsew
rlabel metal1 s 9726 16960 9762 17301 4 vdd
port 515 nsew
rlabel metal1 s 10206 16669 10242 17010 4 vdd
port 515 nsew
rlabel metal1 s 6462 9559 6498 9900 4 vdd
port 515 nsew
rlabel metal1 s 4734 869 4770 1210 4 vdd
port 515 nsew
rlabel metal1 s 4734 8270 4770 8611 4 vdd
port 515 nsew
rlabel metal1 s 222 3239 258 3580 4 vdd
port 515 nsew
rlabel metal1 s 16446 4819 16482 5160 4 vdd
port 515 nsew
rlabel metal1 s 14718 14590 14754 14931 4 vdd
port 515 nsew
rlabel metal1 s 9726 24070 9762 24411 4 vdd
port 515 nsew
rlabel metal1 s 16446 10349 16482 10690 4 vdd
port 515 nsew
rlabel metal1 s 16446 20910 16482 21251 4 vdd
port 515 nsew
rlabel metal1 s 11454 12220 11490 12561 4 vdd
port 515 nsew
rlabel metal1 s 19710 18540 19746 18881 4 vdd
port 515 nsew
rlabel metal1 s 8958 9559 8994 9900 4 vdd
port 515 nsew
rlabel metal1 s 5982 19330 6018 19671 4 vdd
port 515 nsew
rlabel metal1 s 7230 20120 7266 20461 4 vdd
port 515 nsew
rlabel metal1 s 11454 23779 11490 24120 4 vdd
port 515 nsew
rlabel metal1 s 18942 3530 18978 3871 4 vdd
port 515 nsew
rlabel metal1 s 17694 1950 17730 2291 4 vdd
port 515 nsew
rlabel metal1 s 3966 7480 4002 7821 4 vdd
port 515 nsew
rlabel metal1 s 222 5110 258 5451 4 vdd
port 515 nsew
rlabel metal1 s 11454 20910 11490 21251 4 vdd
port 515 nsew
rlabel metal1 s 5982 23280 6018 23621 4 vdd
port 515 nsew
rlabel metal1 s 222 7480 258 7821 4 vdd
port 515 nsew
rlabel metal1 s 13950 19330 13986 19671 4 vdd
port 515 nsew
rlabel metal1 s 5982 13010 6018 13351 4 vdd
port 515 nsew
rlabel metal1 s 18942 22490 18978 22831 4 vdd
port 515 nsew
rlabel metal1 s 2238 19039 2274 19380 4 vdd
port 515 nsew
rlabel metal1 s 17694 4320 17730 4661 4 vdd
port 515 nsew
rlabel metal1 s 7710 8769 7746 9110 4 vdd
port 515 nsew
rlabel metal1 s 9726 7480 9762 7821 4 vdd
port 515 nsew
rlabel metal1 s 17214 9060 17250 9401 4 vdd
port 515 nsew
rlabel metal1 s 10206 19829 10242 20170 4 vdd
port 515 nsew
rlabel metal1 s 12222 7189 12258 7530 4 vdd
port 515 nsew
rlabel metal1 s 1470 11430 1506 11771 4 vdd
port 515 nsew
rlabel metal1 s 10206 12220 10242 12561 4 vdd
port 515 nsew
rlabel metal1 s 17694 8270 17730 8611 4 vdd
port 515 nsew
rlabel metal1 s 3486 15089 3522 15430 4 vdd
port 515 nsew
rlabel metal1 s 18942 5900 18978 6241 4 vdd
port 515 nsew
rlabel metal1 s 19710 23779 19746 24120 4 vdd
port 515 nsew
rlabel metal1 s 12702 1160 12738 1501 4 vdd
port 515 nsew
rlabel metal1 s 1470 19039 1506 19380 4 vdd
port 515 nsew
rlabel metal1 s 5214 21700 5250 22041 4 vdd
port 515 nsew
rlabel metal1 s 18462 5110 18498 5451 4 vdd
port 515 nsew
rlabel metal1 s 8478 13010 8514 13351 4 vdd
port 515 nsew
rlabel metal1 s 3966 14590 4002 14931 4 vdd
port 515 nsew
rlabel metal1 s 15198 7480 15234 7821 4 vdd
port 515 nsew
rlabel metal1 s 2238 15879 2274 16220 4 vdd
port 515 nsew
rlabel metal1 s 12702 5900 12738 6241 4 vdd
port 515 nsew
rlabel metal1 s 12222 15380 12258 15721 4 vdd
port 515 nsew
rlabel metal1 s 5214 4320 5250 4661 4 vdd
port 515 nsew
rlabel metal1 s 16446 11929 16482 12270 4 vdd
port 515 nsew
rlabel metal1 s 9726 3239 9762 3580 4 vdd
port 515 nsew
rlabel metal1 s 10974 4029 11010 4370 4 vdd
port 515 nsew
rlabel metal1 s 12222 1160 12258 1501 4 vdd
port 515 nsew
rlabel metal1 s 12222 7979 12258 8320 4 vdd
port 515 nsew
rlabel metal1 s 19710 13010 19746 13351 4 vdd
port 515 nsew
rlabel metal1 s 14718 12719 14754 13060 4 vdd
port 515 nsew
rlabel metal1 s 10974 1659 11010 2000 4 vdd
port 515 nsew
rlabel metal1 s 10206 11139 10242 11480 4 vdd
port 515 nsew
rlabel metal1 s 13950 12719 13986 13060 4 vdd
port 515 nsew
rlabel metal1 s 17694 1160 17730 1501 4 vdd
port 515 nsew
rlabel metal1 s 2718 11139 2754 11480 4 vdd
port 515 nsew
rlabel metal1 s 12222 18249 12258 18590 4 vdd
port 515 nsew
rlabel metal1 s 222 869 258 1210 4 vdd
port 515 nsew
rlabel metal1 s 4734 14299 4770 14640 4 vdd
port 515 nsew
rlabel metal1 s 9726 19039 9762 19380 4 vdd
port 515 nsew
rlabel metal1 s 4734 16960 4770 17301 4 vdd
port 515 nsew
rlabel metal1 s 17214 20619 17250 20960 4 vdd
port 515 nsew
rlabel metal1 s 8958 21700 8994 22041 4 vdd
port 515 nsew
rlabel metal1 s 10206 1950 10242 2291 4 vdd
port 515 nsew
rlabel metal1 s 14718 20910 14754 21251 4 vdd
port 515 nsew
rlabel metal1 s 16446 20120 16482 20461 4 vdd
port 515 nsew
rlabel metal1 s 16446 22199 16482 22540 4 vdd
port 515 nsew
rlabel metal1 s 6462 4819 6498 5160 4 vdd
port 515 nsew
rlabel metal1 s 222 20120 258 20461 4 vdd
port 515 nsew
rlabel metal1 s 5982 370 6018 711 4 vdd
port 515 nsew
rlabel metal1 s 19710 17750 19746 18091 4 vdd
port 515 nsew
rlabel metal1 s 15198 22989 15234 23330 4 vdd
port 515 nsew
rlabel metal1 s 2238 13010 2274 13351 4 vdd
port 515 nsew
rlabel metal1 s 8478 12220 8514 12561 4 vdd
port 515 nsew
rlabel metal1 s 17214 79 17250 420 4 vdd
port 515 nsew
rlabel metal1 s 4734 8769 4770 9110 4 vdd
port 515 nsew
rlabel metal1 s 4734 13800 4770 14141 4 vdd
port 515 nsew
rlabel metal1 s 17694 18540 17730 18881 4 vdd
port 515 nsew
rlabel metal1 s 222 4819 258 5160 4 vdd
port 515 nsew
rlabel metal1 s 15198 24569 15234 24910 4 vdd
port 515 nsew
rlabel metal1 s 19710 24070 19746 24411 4 vdd
port 515 nsew
rlabel metal1 s 222 6399 258 6740 4 vdd
port 515 nsew
rlabel metal1 s 12222 6399 12258 6740 4 vdd
port 515 nsew
rlabel metal1 s 15198 24070 15234 24411 4 vdd
port 515 nsew
rlabel metal1 s 6462 19829 6498 20170 4 vdd
port 515 nsew
rlabel metal1 s 6462 18540 6498 18881 4 vdd
port 515 nsew
rlabel metal1 s 3966 3530 4002 3871 4 vdd
port 515 nsew
rlabel metal1 s 13470 3239 13506 3580 4 vdd
port 515 nsew
rlabel metal1 s 14718 1950 14754 2291 4 vdd
port 515 nsew
rlabel metal1 s 5982 18540 6018 18881 4 vdd
port 515 nsew
rlabel metal1 s 18942 24070 18978 24411 4 vdd
port 515 nsew
rlabel metal1 s 3966 15380 4002 15721 4 vdd
port 515 nsew
rlabel metal1 s 9726 20619 9762 20960 4 vdd
port 515 nsew
rlabel metal1 s 13950 23280 13986 23621 4 vdd
port 515 nsew
rlabel metal1 s 222 13010 258 13351 4 vdd
port 515 nsew
rlabel metal1 s 222 18540 258 18881 4 vdd
port 515 nsew
rlabel metal1 s 2718 21700 2754 22041 4 vdd
port 515 nsew
rlabel metal1 s 3966 6399 4002 6740 4 vdd
port 515 nsew
rlabel metal1 s 2718 10349 2754 10690 4 vdd
port 515 nsew
rlabel metal1 s 990 19829 1026 20170 4 vdd
port 515 nsew
rlabel metal1 s 990 11430 1026 11771 4 vdd
port 515 nsew
rlabel metal1 s 15966 2449 16002 2790 4 vdd
port 515 nsew
rlabel metal1 s 17694 2740 17730 3081 4 vdd
port 515 nsew
rlabel metal1 s 10206 21409 10242 21750 4 vdd
port 515 nsew
rlabel metal1 s 1470 16170 1506 16511 4 vdd
port 515 nsew
rlabel metal1 s 2238 79 2274 420 4 vdd
port 515 nsew
rlabel metal1 s 17694 10640 17730 10981 4 vdd
port 515 nsew
rlabel metal1 s 5982 19829 6018 20170 4 vdd
port 515 nsew
rlabel metal1 s 2238 16170 2274 16511 4 vdd
port 515 nsew
rlabel metal1 s 19710 13800 19746 14141 4 vdd
port 515 nsew
rlabel metal1 s 7710 14590 7746 14931 4 vdd
port 515 nsew
rlabel metal1 s 14718 7480 14754 7821 4 vdd
port 515 nsew
rlabel metal1 s 2238 4029 2274 4370 4 vdd
port 515 nsew
rlabel metal1 s 9726 8769 9762 9110 4 vdd
port 515 nsew
rlabel metal1 s 18942 15380 18978 15721 4 vdd
port 515 nsew
rlabel metal1 s 10974 20619 11010 20960 4 vdd
port 515 nsew
rlabel metal1 s 1470 12719 1506 13060 4 vdd
port 515 nsew
rlabel metal1 s 18462 20910 18498 21251 4 vdd
port 515 nsew
rlabel metal1 s 6462 23280 6498 23621 4 vdd
port 515 nsew
rlabel metal1 s 19710 23280 19746 23621 4 vdd
port 515 nsew
rlabel metal1 s 15198 1160 15234 1501 4 vdd
port 515 nsew
rlabel metal1 s 13470 14299 13506 14640 4 vdd
port 515 nsew
rlabel metal1 s 18942 6690 18978 7031 4 vdd
port 515 nsew
rlabel metal1 s 17214 20910 17250 21251 4 vdd
port 515 nsew
rlabel metal1 s 17214 15879 17250 16220 4 vdd
port 515 nsew
rlabel metal1 s 15198 10640 15234 10981 4 vdd
port 515 nsew
rlabel metal1 s 15966 14299 16002 14640 4 vdd
port 515 nsew
rlabel metal1 s 7230 7480 7266 7821 4 vdd
port 515 nsew
rlabel metal1 s 18462 5900 18498 6241 4 vdd
port 515 nsew
rlabel metal1 s 5982 7480 6018 7821 4 vdd
port 515 nsew
rlabel metal1 s 1470 20910 1506 21251 4 vdd
port 515 nsew
rlabel metal1 s 13470 5900 13506 6241 4 vdd
port 515 nsew
rlabel metal1 s 17214 10640 17250 10981 4 vdd
port 515 nsew
rlabel metal1 s 10206 24569 10242 24910 4 vdd
port 515 nsew
rlabel metal1 s 13950 18249 13986 18590 4 vdd
port 515 nsew
rlabel metal1 s 11454 20120 11490 20461 4 vdd
port 515 nsew
rlabel metal1 s 8478 14590 8514 14931 4 vdd
port 515 nsew
rlabel metal1 s 17214 6399 17250 6740 4 vdd
port 515 nsew
rlabel metal1 s 222 16170 258 16511 4 vdd
port 515 nsew
rlabel metal1 s 19710 9060 19746 9401 4 vdd
port 515 nsew
rlabel metal1 s 5214 15879 5250 16220 4 vdd
port 515 nsew
rlabel metal1 s 7710 20619 7746 20960 4 vdd
port 515 nsew
rlabel metal1 s 8958 869 8994 1210 4 vdd
port 515 nsew
rlabel metal1 s 990 19039 1026 19380 4 vdd
port 515 nsew
rlabel metal1 s 16446 370 16482 711 4 vdd
port 515 nsew
rlabel metal1 s 13950 5900 13986 6241 4 vdd
port 515 nsew
rlabel metal1 s 15198 13509 15234 13850 4 vdd
port 515 nsew
rlabel metal1 s 15966 23280 16002 23621 4 vdd
port 515 nsew
rlabel metal1 s 990 4819 1026 5160 4 vdd
port 515 nsew
rlabel metal1 s 7710 24070 7746 24411 4 vdd
port 515 nsew
rlabel metal1 s 5214 10349 5250 10690 4 vdd
port 515 nsew
rlabel metal1 s 11454 79 11490 420 4 vdd
port 515 nsew
rlabel metal1 s 15198 2740 15234 3081 4 vdd
port 515 nsew
rlabel metal1 s 17214 22199 17250 22540 4 vdd
port 515 nsew
rlabel metal1 s 12222 15089 12258 15430 4 vdd
port 515 nsew
rlabel metal1 s 222 79 258 420 4 vdd
port 515 nsew
rlabel metal1 s 13950 5110 13986 5451 4 vdd
port 515 nsew
rlabel metal1 s 4734 24070 4770 24411 4 vdd
port 515 nsew
rlabel metal1 s 222 17750 258 18091 4 vdd
port 515 nsew
rlabel metal1 s 15966 6690 16002 7031 4 vdd
port 515 nsew
rlabel metal1 s 3486 19330 3522 19671 4 vdd
port 515 nsew
rlabel metal1 s 10206 2740 10242 3081 4 vdd
port 515 nsew
rlabel metal1 s 222 24070 258 24411 4 vdd
port 515 nsew
rlabel metal1 s 17214 1659 17250 2000 4 vdd
port 515 nsew
rlabel metal1 s 4734 22199 4770 22540 4 vdd
port 515 nsew
rlabel metal1 s 3966 18540 4002 18881 4 vdd
port 515 nsew
rlabel metal1 s 2718 4819 2754 5160 4 vdd
port 515 nsew
rlabel metal1 s 13950 5609 13986 5950 4 vdd
port 515 nsew
rlabel metal1 s 19710 11139 19746 11480 4 vdd
port 515 nsew
rlabel metal1 s 18942 18540 18978 18881 4 vdd
port 515 nsew
rlabel metal1 s 18462 12719 18498 13060 4 vdd
port 515 nsew
rlabel metal1 s 15966 11139 16002 11480 4 vdd
port 515 nsew
rlabel metal1 s 19710 22989 19746 23330 4 vdd
port 515 nsew
rlabel metal1 s 5214 12719 5250 13060 4 vdd
port 515 nsew
rlabel metal1 s 2238 22199 2274 22540 4 vdd
port 515 nsew
rlabel metal1 s 3966 79 4002 420 4 vdd
port 515 nsew
rlabel metal1 s 4734 15089 4770 15430 4 vdd
port 515 nsew
rlabel metal1 s 13950 22199 13986 22540 4 vdd
port 515 nsew
rlabel metal1 s 3966 19039 4002 19380 4 vdd
port 515 nsew
rlabel metal1 s 990 3530 1026 3871 4 vdd
port 515 nsew
rlabel metal1 s 3486 370 3522 711 4 vdd
port 515 nsew
rlabel metal1 s 13950 4029 13986 4370 4 vdd
port 515 nsew
rlabel metal1 s 990 22989 1026 23330 4 vdd
port 515 nsew
rlabel metal1 s 5982 9060 6018 9401 4 vdd
port 515 nsew
rlabel metal1 s 4734 5900 4770 6241 4 vdd
port 515 nsew
rlabel metal1 s 15198 21700 15234 22041 4 vdd
port 515 nsew
rlabel metal1 s 2238 18249 2274 18590 4 vdd
port 515 nsew
rlabel metal1 s 4734 21409 4770 21750 4 vdd
port 515 nsew
rlabel metal1 s 7230 24070 7266 24411 4 vdd
port 515 nsew
rlabel metal1 s 17214 8270 17250 8611 4 vdd
port 515 nsew
rlabel metal1 s 5214 17459 5250 17800 4 vdd
port 515 nsew
rlabel metal1 s 2718 15089 2754 15430 4 vdd
port 515 nsew
rlabel metal1 s 2238 5609 2274 5950 4 vdd
port 515 nsew
rlabel metal1 s 1470 21409 1506 21750 4 vdd
port 515 nsew
rlabel metal1 s 18462 1160 18498 1501 4 vdd
port 515 nsew
rlabel metal1 s 5214 16170 5250 16511 4 vdd
port 515 nsew
rlabel metal1 s 13470 20120 13506 20461 4 vdd
port 515 nsew
rlabel metal1 s 2718 3530 2754 3871 4 vdd
port 515 nsew
rlabel metal1 s 16446 6690 16482 7031 4 vdd
port 515 nsew
rlabel metal1 s 12702 20910 12738 21251 4 vdd
port 515 nsew
rlabel metal1 s 17694 5609 17730 5950 4 vdd
port 515 nsew
rlabel metal1 s 1470 1160 1506 1501 4 vdd
port 515 nsew
rlabel metal1 s 1470 12220 1506 12561 4 vdd
port 515 nsew
rlabel metal1 s 990 5110 1026 5451 4 vdd
port 515 nsew
rlabel metal1 s 13470 16960 13506 17301 4 vdd
port 515 nsew
rlabel metal1 s 2238 1659 2274 2000 4 vdd
port 515 nsew
rlabel metal1 s 13470 16170 13506 16511 4 vdd
port 515 nsew
rlabel metal1 s 6462 5110 6498 5451 4 vdd
port 515 nsew
rlabel metal1 s 17694 1659 17730 2000 4 vdd
port 515 nsew
rlabel metal1 s 2238 17459 2274 17800 4 vdd
port 515 nsew
rlabel metal1 s 8958 11139 8994 11480 4 vdd
port 515 nsew
rlabel metal1 s 10974 7189 11010 7530 4 vdd
port 515 nsew
rlabel metal1 s 1470 22989 1506 23330 4 vdd
port 515 nsew
rlabel metal1 s 18462 10640 18498 10981 4 vdd
port 515 nsew
rlabel metal1 s 3966 19829 4002 20170 4 vdd
port 515 nsew
rlabel metal1 s 5982 9559 6018 9900 4 vdd
port 515 nsew
rlabel metal1 s 18462 22989 18498 23330 4 vdd
port 515 nsew
rlabel metal1 s 13950 17750 13986 18091 4 vdd
port 515 nsew
rlabel metal1 s 13470 24860 13506 25201 4 vdd
port 515 nsew
rlabel metal1 s 12702 9060 12738 9401 4 vdd
port 515 nsew
rlabel metal1 s 15966 22989 16002 23330 4 vdd
port 515 nsew
rlabel metal1 s 7710 24569 7746 24910 4 vdd
port 515 nsew
rlabel metal1 s 2238 8270 2274 8611 4 vdd
port 515 nsew
rlabel metal1 s 222 8270 258 8611 4 vdd
port 515 nsew
rlabel metal1 s 16446 12719 16482 13060 4 vdd
port 515 nsew
rlabel metal1 s 13470 24569 13506 24910 4 vdd
port 515 nsew
rlabel metal1 s 7230 17459 7266 17800 4 vdd
port 515 nsew
rlabel metal1 s 7710 1659 7746 2000 4 vdd
port 515 nsew
rlabel metal1 s 8958 5609 8994 5950 4 vdd
port 515 nsew
rlabel metal1 s 15198 8769 15234 9110 4 vdd
port 515 nsew
rlabel metal1 s 9726 13800 9762 14141 4 vdd
port 515 nsew
rlabel metal1 s 12222 22490 12258 22831 4 vdd
port 515 nsew
rlabel metal1 s 8958 13010 8994 13351 4 vdd
port 515 nsew
rlabel metal1 s 13470 22199 13506 22540 4 vdd
port 515 nsew
rlabel metal1 s 15198 15879 15234 16220 4 vdd
port 515 nsew
rlabel metal1 s 18462 3530 18498 3871 4 vdd
port 515 nsew
rlabel metal1 s 10974 8769 11010 9110 4 vdd
port 515 nsew
rlabel metal1 s 2238 12719 2274 13060 4 vdd
port 515 nsew
rlabel metal1 s 222 1950 258 2291 4 vdd
port 515 nsew
rlabel metal1 s 7230 1659 7266 2000 4 vdd
port 515 nsew
rlabel metal1 s 3966 2449 4002 2790 4 vdd
port 515 nsew
rlabel metal1 s 12702 18249 12738 18590 4 vdd
port 515 nsew
rlabel metal1 s 1470 19829 1506 20170 4 vdd
port 515 nsew
rlabel metal1 s 17214 16960 17250 17301 4 vdd
port 515 nsew
rlabel metal1 s 8958 4320 8994 4661 4 vdd
port 515 nsew
rlabel metal1 s 14718 869 14754 1210 4 vdd
port 515 nsew
rlabel metal1 s 6462 79 6498 420 4 vdd
port 515 nsew
rlabel metal1 s 15966 19829 16002 20170 4 vdd
port 515 nsew
rlabel metal1 s 4734 20910 4770 21251 4 vdd
port 515 nsew
rlabel metal1 s 3486 16960 3522 17301 4 vdd
port 515 nsew
rlabel metal1 s 15198 4819 15234 5160 4 vdd
port 515 nsew
rlabel metal1 s 12222 13800 12258 14141 4 vdd
port 515 nsew
rlabel metal1 s 6462 12719 6498 13060 4 vdd
port 515 nsew
rlabel metal1 s 3486 3530 3522 3871 4 vdd
port 515 nsew
rlabel metal1 s 18942 16170 18978 16511 4 vdd
port 515 nsew
rlabel metal1 s 7710 1950 7746 2291 4 vdd
port 515 nsew
rlabel metal1 s 13470 24070 13506 24411 4 vdd
port 515 nsew
rlabel metal1 s 4734 5609 4770 5950 4 vdd
port 515 nsew
rlabel metal1 s 17214 13010 17250 13351 4 vdd
port 515 nsew
rlabel metal1 s 10206 18249 10242 18590 4 vdd
port 515 nsew
rlabel metal1 s 11454 1659 11490 2000 4 vdd
port 515 nsew
rlabel metal1 s 11454 21700 11490 22041 4 vdd
port 515 nsew
rlabel metal1 s 3966 9850 4002 10191 4 vdd
port 515 nsew
rlabel metal1 s 5982 22989 6018 23330 4 vdd
port 515 nsew
rlabel metal1 s 7710 5110 7746 5451 4 vdd
port 515 nsew
rlabel metal1 s 3966 21700 4002 22041 4 vdd
port 515 nsew
rlabel metal1 s 17214 22490 17250 22831 4 vdd
port 515 nsew
rlabel metal1 s 12702 6690 12738 7031 4 vdd
port 515 nsew
rlabel metal1 s 990 13509 1026 13850 4 vdd
port 515 nsew
rlabel metal1 s 16446 1659 16482 2000 4 vdd
port 515 nsew
rlabel metal1 s 15966 24070 16002 24411 4 vdd
port 515 nsew
rlabel metal1 s 18462 4029 18498 4370 4 vdd
port 515 nsew
rlabel metal1 s 8478 15089 8514 15430 4 vdd
port 515 nsew
rlabel metal1 s 7710 7480 7746 7821 4 vdd
port 515 nsew
rlabel metal1 s 990 8769 1026 9110 4 vdd
port 515 nsew
rlabel metal1 s 7230 4819 7266 5160 4 vdd
port 515 nsew
rlabel metal1 s 222 15089 258 15430 4 vdd
port 515 nsew
rlabel metal1 s 9726 15879 9762 16220 4 vdd
port 515 nsew
rlabel metal1 s 4734 1160 4770 1501 4 vdd
port 515 nsew
rlabel metal1 s 8958 9850 8994 10191 4 vdd
port 515 nsew
rlabel metal1 s 6462 14590 6498 14931 4 vdd
port 515 nsew
rlabel metal1 s 8478 20910 8514 21251 4 vdd
port 515 nsew
rlabel metal1 s 17214 16669 17250 17010 4 vdd
port 515 nsew
rlabel metal1 s 12222 21409 12258 21750 4 vdd
port 515 nsew
rlabel metal1 s 8478 15879 8514 16220 4 vdd
port 515 nsew
rlabel metal1 s 2238 24569 2274 24910 4 vdd
port 515 nsew
rlabel metal1 s 8958 4029 8994 4370 4 vdd
port 515 nsew
rlabel metal1 s 9726 869 9762 1210 4 vdd
port 515 nsew
rlabel metal1 s 11454 22989 11490 23330 4 vdd
port 515 nsew
rlabel metal1 s 16446 14299 16482 14640 4 vdd
port 515 nsew
rlabel metal1 s 12222 22989 12258 23330 4 vdd
port 515 nsew
rlabel metal1 s 7710 13800 7746 14141 4 vdd
port 515 nsew
rlabel metal1 s 1470 22490 1506 22831 4 vdd
port 515 nsew
rlabel metal1 s 10206 24070 10242 24411 4 vdd
port 515 nsew
rlabel metal1 s 8958 23779 8994 24120 4 vdd
port 515 nsew
rlabel metal1 s 6462 6399 6498 6740 4 vdd
port 515 nsew
rlabel metal1 s 10206 4819 10242 5160 4 vdd
port 515 nsew
rlabel metal1 s 5214 7189 5250 7530 4 vdd
port 515 nsew
rlabel metal1 s 9726 1160 9762 1501 4 vdd
port 515 nsew
rlabel metal1 s 17214 1160 17250 1501 4 vdd
port 515 nsew
rlabel metal1 s 17214 370 17250 711 4 vdd
port 515 nsew
rlabel metal1 s 14718 17750 14754 18091 4 vdd
port 515 nsew
rlabel metal1 s 3486 1659 3522 2000 4 vdd
port 515 nsew
rlabel metal1 s 2718 15879 2754 16220 4 vdd
port 515 nsew
rlabel metal1 s 13470 9060 13506 9401 4 vdd
port 515 nsew
rlabel metal1 s 9726 5900 9762 6241 4 vdd
port 515 nsew
rlabel metal1 s 13950 4320 13986 4661 4 vdd
port 515 nsew
rlabel metal1 s 13950 24860 13986 25201 4 vdd
port 515 nsew
rlabel metal1 s 3486 17459 3522 17800 4 vdd
port 515 nsew
rlabel metal1 s 16446 5110 16482 5451 4 vdd
port 515 nsew
rlabel metal1 s 14718 24860 14754 25201 4 vdd
port 515 nsew
rlabel metal1 s 9726 14590 9762 14931 4 vdd
port 515 nsew
rlabel metal1 s 13950 15089 13986 15430 4 vdd
port 515 nsew
rlabel metal1 s 990 24070 1026 24411 4 vdd
port 515 nsew
rlabel metal1 s 5982 21700 6018 22041 4 vdd
port 515 nsew
rlabel metal1 s 12702 24860 12738 25201 4 vdd
port 515 nsew
rlabel metal1 s 2718 5110 2754 5451 4 vdd
port 515 nsew
rlabel metal1 s 15966 13800 16002 14141 4 vdd
port 515 nsew
rlabel metal1 s 2718 13509 2754 13850 4 vdd
port 515 nsew
rlabel metal1 s 19710 869 19746 1210 4 vdd
port 515 nsew
rlabel metal1 s 9726 20910 9762 21251 4 vdd
port 515 nsew
rlabel metal1 s 222 5900 258 6241 4 vdd
port 515 nsew
rlabel metal1 s 5214 15380 5250 15721 4 vdd
port 515 nsew
rlabel metal1 s 2238 2740 2274 3081 4 vdd
port 515 nsew
rlabel metal1 s 17694 12220 17730 12561 4 vdd
port 515 nsew
rlabel metal1 s 12702 23779 12738 24120 4 vdd
port 515 nsew
rlabel metal1 s 4734 9060 4770 9401 4 vdd
port 515 nsew
rlabel metal1 s 12222 9559 12258 9900 4 vdd
port 515 nsew
rlabel metal1 s 8958 21409 8994 21750 4 vdd
port 515 nsew
rlabel metal1 s 8478 3239 8514 3580 4 vdd
port 515 nsew
rlabel metal1 s 990 11139 1026 11480 4 vdd
port 515 nsew
rlabel metal1 s 12702 79 12738 420 4 vdd
port 515 nsew
rlabel metal1 s 13470 7189 13506 7530 4 vdd
port 515 nsew
rlabel metal1 s 5214 10640 5250 10981 4 vdd
port 515 nsew
rlabel metal1 s 14718 11430 14754 11771 4 vdd
port 515 nsew
rlabel metal1 s 8478 16960 8514 17301 4 vdd
port 515 nsew
rlabel metal1 s 8478 23779 8514 24120 4 vdd
port 515 nsew
rlabel metal1 s 3966 12719 4002 13060 4 vdd
port 515 nsew
rlabel metal1 s 7710 19829 7746 20170 4 vdd
port 515 nsew
rlabel metal1 s 3966 17459 4002 17800 4 vdd
port 515 nsew
rlabel metal1 s 4734 17459 4770 17800 4 vdd
port 515 nsew
rlabel metal1 s 13470 15380 13506 15721 4 vdd
port 515 nsew
rlabel metal1 s 5982 17459 6018 17800 4 vdd
port 515 nsew
rlabel metal1 s 16446 3239 16482 3580 4 vdd
port 515 nsew
rlabel metal1 s 7710 22199 7746 22540 4 vdd
port 515 nsew
rlabel metal1 s 1470 7480 1506 7821 4 vdd
port 515 nsew
rlabel metal1 s 5214 8270 5250 8611 4 vdd
port 515 nsew
rlabel metal1 s 7230 4320 7266 4661 4 vdd
port 515 nsew
rlabel metal1 s 15966 13010 16002 13351 4 vdd
port 515 nsew
rlabel metal1 s 990 13800 1026 14141 4 vdd
port 515 nsew
rlabel metal1 s 19710 2740 19746 3081 4 vdd
port 515 nsew
rlabel metal1 s 1470 1950 1506 2291 4 vdd
port 515 nsew
rlabel metal1 s 13950 4819 13986 5160 4 vdd
port 515 nsew
rlabel metal1 s 15966 6399 16002 6740 4 vdd
port 515 nsew
rlabel metal1 s 19710 12220 19746 12561 4 vdd
port 515 nsew
rlabel metal1 s 12702 8270 12738 8611 4 vdd
port 515 nsew
rlabel metal1 s 8478 17459 8514 17800 4 vdd
port 515 nsew
rlabel metal1 s 13470 18249 13506 18590 4 vdd
port 515 nsew
rlabel metal1 s 14718 79 14754 420 4 vdd
port 515 nsew
rlabel metal1 s 18462 20619 18498 20960 4 vdd
port 515 nsew
rlabel metal1 s 18462 14590 18498 14931 4 vdd
port 515 nsew
rlabel metal1 s 1470 17750 1506 18091 4 vdd
port 515 nsew
rlabel metal1 s 7230 12220 7266 12561 4 vdd
port 515 nsew
rlabel metal1 s 2718 16170 2754 16511 4 vdd
port 515 nsew
rlabel metal1 s 14718 16669 14754 17010 4 vdd
port 515 nsew
rlabel metal1 s 2718 19039 2754 19380 4 vdd
port 515 nsew
rlabel metal1 s 18942 8270 18978 8611 4 vdd
port 515 nsew
rlabel metal1 s 10206 5900 10242 6241 4 vdd
port 515 nsew
rlabel metal1 s 3966 5110 4002 5451 4 vdd
port 515 nsew
rlabel metal1 s 4734 4029 4770 4370 4 vdd
port 515 nsew
rlabel metal1 s 8958 1160 8994 1501 4 vdd
port 515 nsew
rlabel metal1 s 5214 19039 5250 19380 4 vdd
port 515 nsew
rlabel metal1 s 11454 16669 11490 17010 4 vdd
port 515 nsew
rlabel metal1 s 14718 14299 14754 14640 4 vdd
port 515 nsew
rlabel metal1 s 2238 19829 2274 20170 4 vdd
port 515 nsew
rlabel metal1 s 3486 24569 3522 24910 4 vdd
port 515 nsew
rlabel metal1 s 3486 23280 3522 23621 4 vdd
port 515 nsew
rlabel metal1 s 2718 3239 2754 3580 4 vdd
port 515 nsew
rlabel metal1 s 5982 869 6018 1210 4 vdd
port 515 nsew
rlabel metal1 s 10974 11430 11010 11771 4 vdd
port 515 nsew
rlabel metal1 s 19710 4029 19746 4370 4 vdd
port 515 nsew
rlabel metal1 s 15966 1160 16002 1501 4 vdd
port 515 nsew
rlabel metal1 s 10974 18249 11010 18590 4 vdd
port 515 nsew
rlabel metal1 s 17214 5110 17250 5451 4 vdd
port 515 nsew
rlabel metal1 s 222 24569 258 24910 4 vdd
port 515 nsew
rlabel metal1 s 5214 22490 5250 22831 4 vdd
port 515 nsew
rlabel metal1 s 7230 869 7266 1210 4 vdd
port 515 nsew
rlabel metal1 s 3486 21409 3522 21750 4 vdd
port 515 nsew
rlabel metal1 s 7710 12220 7746 12561 4 vdd
port 515 nsew
rlabel metal1 s 17214 4819 17250 5160 4 vdd
port 515 nsew
rlabel metal1 s 3966 370 4002 711 4 vdd
port 515 nsew
rlabel metal1 s 4734 23779 4770 24120 4 vdd
port 515 nsew
rlabel metal1 s 7710 24860 7746 25201 4 vdd
port 515 nsew
rlabel metal1 s 17694 14299 17730 14640 4 vdd
port 515 nsew
rlabel metal1 s 14718 3239 14754 3580 4 vdd
port 515 nsew
rlabel metal1 s 3486 12719 3522 13060 4 vdd
port 515 nsew
rlabel metal1 s 19710 3530 19746 3871 4 vdd
port 515 nsew
rlabel metal1 s 17214 4320 17250 4661 4 vdd
port 515 nsew
rlabel metal1 s 17694 4029 17730 4370 4 vdd
port 515 nsew
rlabel metal1 s 19710 20120 19746 20461 4 vdd
port 515 nsew
rlabel metal1 s 5214 9850 5250 10191 4 vdd
port 515 nsew
rlabel metal1 s 10974 22199 11010 22540 4 vdd
port 515 nsew
rlabel metal1 s 1470 4819 1506 5160 4 vdd
port 515 nsew
rlabel metal1 s 13470 17459 13506 17800 4 vdd
port 515 nsew
rlabel metal1 s 17694 15879 17730 16220 4 vdd
port 515 nsew
rlabel metal1 s 13470 9850 13506 10191 4 vdd
port 515 nsew
rlabel metal1 s 14718 3530 14754 3871 4 vdd
port 515 nsew
rlabel metal1 s 3486 20910 3522 21251 4 vdd
port 515 nsew
rlabel metal1 s 8478 1160 8514 1501 4 vdd
port 515 nsew
rlabel metal1 s 12222 23779 12258 24120 4 vdd
port 515 nsew
rlabel metal1 s 2718 869 2754 1210 4 vdd
port 515 nsew
rlabel metal1 s 14718 15380 14754 15721 4 vdd
port 515 nsew
rlabel metal1 s 17694 11929 17730 12270 4 vdd
port 515 nsew
rlabel metal1 s 15966 9559 16002 9900 4 vdd
port 515 nsew
rlabel metal1 s 7230 8270 7266 8611 4 vdd
port 515 nsew
rlabel metal1 s 13470 1659 13506 2000 4 vdd
port 515 nsew
rlabel metal1 s 6462 3239 6498 3580 4 vdd
port 515 nsew
rlabel metal1 s 19710 1659 19746 2000 4 vdd
port 515 nsew
rlabel metal1 s 2238 12220 2274 12561 4 vdd
port 515 nsew
rlabel metal1 s 19710 4320 19746 4661 4 vdd
port 515 nsew
rlabel metal1 s 990 6399 1026 6740 4 vdd
port 515 nsew
rlabel metal1 s 19710 16170 19746 16511 4 vdd
port 515 nsew
rlabel metal1 s 13950 2449 13986 2790 4 vdd
port 515 nsew
rlabel metal1 s 17694 22199 17730 22540 4 vdd
port 515 nsew
rlabel metal1 s 17694 23280 17730 23621 4 vdd
port 515 nsew
rlabel metal1 s 2718 19829 2754 20170 4 vdd
port 515 nsew
rlabel metal1 s 2718 11929 2754 12270 4 vdd
port 515 nsew
rlabel metal1 s 14718 8769 14754 9110 4 vdd
port 515 nsew
rlabel metal1 s 15198 9060 15234 9401 4 vdd
port 515 nsew
rlabel metal1 s 6462 11430 6498 11771 4 vdd
port 515 nsew
rlabel metal1 s 7230 21700 7266 22041 4 vdd
port 515 nsew
rlabel metal1 s 5214 20120 5250 20461 4 vdd
port 515 nsew
rlabel metal1 s 1470 5609 1506 5950 4 vdd
port 515 nsew
rlabel metal1 s 8478 24569 8514 24910 4 vdd
port 515 nsew
rlabel metal1 s 11454 15089 11490 15430 4 vdd
port 515 nsew
rlabel metal1 s 3486 10640 3522 10981 4 vdd
port 515 nsew
rlabel metal1 s 2238 18540 2274 18881 4 vdd
port 515 nsew
rlabel metal1 s 7230 15879 7266 16220 4 vdd
port 515 nsew
rlabel metal1 s 7230 1950 7266 2291 4 vdd
port 515 nsew
rlabel metal1 s 6462 2449 6498 2790 4 vdd
port 515 nsew
rlabel metal1 s 19710 19039 19746 19380 4 vdd
port 515 nsew
rlabel metal1 s 2718 8769 2754 9110 4 vdd
port 515 nsew
rlabel metal1 s 2238 15380 2274 15721 4 vdd
port 515 nsew
rlabel metal1 s 16446 9060 16482 9401 4 vdd
port 515 nsew
rlabel metal1 s 9726 18540 9762 18881 4 vdd
port 515 nsew
rlabel metal1 s 990 17750 1026 18091 4 vdd
port 515 nsew
rlabel metal1 s 990 20619 1026 20960 4 vdd
port 515 nsew
rlabel metal1 s 12702 23280 12738 23621 4 vdd
port 515 nsew
rlabel metal1 s 1470 9559 1506 9900 4 vdd
port 515 nsew
rlabel metal1 s 9726 2740 9762 3081 4 vdd
port 515 nsew
rlabel metal1 s 15198 14590 15234 14931 4 vdd
port 515 nsew
rlabel metal1 s 10974 15380 11010 15721 4 vdd
port 515 nsew
rlabel metal1 s 8478 22490 8514 22831 4 vdd
port 515 nsew
rlabel metal1 s 13470 2449 13506 2790 4 vdd
port 515 nsew
rlabel metal1 s 13950 14299 13986 14640 4 vdd
port 515 nsew
rlabel metal1 s 3486 14299 3522 14640 4 vdd
port 515 nsew
rlabel metal1 s 12702 7189 12738 7530 4 vdd
port 515 nsew
rlabel metal1 s 8478 10349 8514 10690 4 vdd
port 515 nsew
rlabel metal1 s 17694 12719 17730 13060 4 vdd
port 515 nsew
rlabel metal1 s 9726 22199 9762 22540 4 vdd
port 515 nsew
rlabel metal1 s 9726 21409 9762 21750 4 vdd
port 515 nsew
rlabel metal1 s 19710 6690 19746 7031 4 vdd
port 515 nsew
rlabel metal1 s 5982 1659 6018 2000 4 vdd
port 515 nsew
rlabel metal1 s 15966 7480 16002 7821 4 vdd
port 515 nsew
rlabel metal1 s 12702 370 12738 711 4 vdd
port 515 nsew
rlabel metal1 s 5214 17750 5250 18091 4 vdd
port 515 nsew
rlabel metal1 s 17694 13010 17730 13351 4 vdd
port 515 nsew
rlabel metal1 s 9726 10640 9762 10981 4 vdd
port 515 nsew
rlabel metal1 s 10974 18540 11010 18881 4 vdd
port 515 nsew
rlabel metal1 s 222 17459 258 17800 4 vdd
port 515 nsew
rlabel metal1 s 18942 20910 18978 21251 4 vdd
port 515 nsew
rlabel metal1 s 2718 1950 2754 2291 4 vdd
port 515 nsew
rlabel metal1 s 10974 3239 11010 3580 4 vdd
port 515 nsew
rlabel metal1 s 16446 16669 16482 17010 4 vdd
port 515 nsew
rlabel metal1 s 17694 24070 17730 24411 4 vdd
port 515 nsew
rlabel metal1 s 3966 13509 4002 13850 4 vdd
port 515 nsew
rlabel metal1 s 13950 13509 13986 13850 4 vdd
port 515 nsew
rlabel metal1 s 17694 20619 17730 20960 4 vdd
port 515 nsew
rlabel metal1 s 1470 23280 1506 23621 4 vdd
port 515 nsew
rlabel metal1 s 3966 20120 4002 20461 4 vdd
port 515 nsew
rlabel metal1 s 222 10640 258 10981 4 vdd
port 515 nsew
rlabel metal1 s 5982 4029 6018 4370 4 vdd
port 515 nsew
rlabel metal1 s 8478 9060 8514 9401 4 vdd
port 515 nsew
rlabel metal1 s 14718 23779 14754 24120 4 vdd
port 515 nsew
rlabel metal1 s 15198 8270 15234 8611 4 vdd
port 515 nsew
rlabel metal1 s 2718 20910 2754 21251 4 vdd
port 515 nsew
rlabel metal1 s 5214 22199 5250 22540 4 vdd
port 515 nsew
rlabel metal1 s 2238 11929 2274 12270 4 vdd
port 515 nsew
rlabel metal1 s 222 7189 258 7530 4 vdd
port 515 nsew
rlabel metal1 s 10974 5900 11010 6241 4 vdd
port 515 nsew
rlabel metal1 s 6462 15380 6498 15721 4 vdd
port 515 nsew
rlabel metal1 s 18462 2740 18498 3081 4 vdd
port 515 nsew
rlabel metal1 s 12222 15879 12258 16220 4 vdd
port 515 nsew
rlabel metal1 s 16446 24860 16482 25201 4 vdd
port 515 nsew
rlabel metal1 s 16446 18249 16482 18590 4 vdd
port 515 nsew
rlabel metal1 s 2718 17750 2754 18091 4 vdd
port 515 nsew
rlabel metal1 s 18942 4819 18978 5160 4 vdd
port 515 nsew
rlabel metal1 s 16446 15089 16482 15430 4 vdd
port 515 nsew
rlabel metal1 s 19710 79 19746 420 4 vdd
port 515 nsew
rlabel metal1 s 16446 19829 16482 20170 4 vdd
port 515 nsew
rlabel metal1 s 5214 19330 5250 19671 4 vdd
port 515 nsew
rlabel metal1 s 9726 6690 9762 7031 4 vdd
port 515 nsew
rlabel metal1 s 15966 15879 16002 16220 4 vdd
port 515 nsew
rlabel metal1 s 3966 15879 4002 16220 4 vdd
port 515 nsew
rlabel metal1 s 3966 2740 4002 3081 4 vdd
port 515 nsew
rlabel metal1 s 12702 24569 12738 24910 4 vdd
port 515 nsew
rlabel metal1 s 2238 7189 2274 7530 4 vdd
port 515 nsew
rlabel metal1 s 6462 5609 6498 5950 4 vdd
port 515 nsew
rlabel metal2 s 14682 6265 14790 6375 4 gnd
port 517 nsew
rlabel metal2 s 17658 17325 17766 17435 4 gnd
port 517 nsew
rlabel metal2 s 3930 20485 4038 20595 4 gnd
port 517 nsew
rlabel metal2 s 12666 5255 12774 5331 4 gnd
port 517 nsew
rlabel metal2 s 12666 12365 12774 12441 4 gnd
port 517 nsew
rlabel metal2 s 6426 7845 6534 7955 4 gnd
port 517 nsew
rlabel metal2 s 186 989 294 1065 4 gnd
port 517 nsew
rlabel metal2 s 3930 24689 4038 24765 4 gnd
port 517 nsew
rlabel metal2 s 6426 21275 6534 21385 4 gnd
port 517 nsew
rlabel metal2 s 2202 17105 2310 17181 4 gnd
port 517 nsew
rlabel metal2 s 5178 22635 5286 22711 4 gnd
port 517 nsew
rlabel metal2 s 15162 12839 15270 12915 4 gnd
port 517 nsew
rlabel metal2 s 6426 17105 6534 17181 4 gnd
port 517 nsew
rlabel metal2 s 3930 15209 4038 15285 4 gnd
port 517 nsew
rlabel metal2 s 12666 18369 12774 18445 4 gnd
port 517 nsew
rlabel metal2 s 12666 18905 12774 19015 4 gnd
port 517 nsew
rlabel metal2 s 17178 12585 17286 12695 4 gnd
port 517 nsew
rlabel metal2 s 17178 12839 17286 12915 4 gnd
port 517 nsew
rlabel metal2 s 4698 11259 4806 11335 4 gnd
port 517 nsew
rlabel metal2 s 186 22635 294 22711 4 gnd
port 517 nsew
rlabel metal2 s 16410 20485 16518 20595 4 gnd
port 517 nsew
rlabel metal2 s 5946 15209 6054 15285 4 gnd
port 517 nsew
rlabel metal2 s 954 7309 1062 7385 4 gnd
port 517 nsew
rlabel metal2 s 186 22855 294 22965 4 gnd
port 517 nsew
rlabel metal2 s 5946 5255 6054 5331 4 gnd
port 517 nsew
rlabel metal2 s 7674 18905 7782 19015 4 gnd
port 517 nsew
rlabel metal2 s 7194 12049 7302 12125 4 gnd
port 517 nsew
rlabel metal2 s 15930 19695 16038 19805 4 gnd
port 517 nsew
rlabel metal2 s 7194 21055 7302 21131 4 gnd
port 517 nsew
rlabel metal2 s 4698 12365 4806 12441 4 gnd
port 517 nsew
rlabel metal2 s 4698 14165 4806 14275 4 gnd
port 517 nsew
rlabel metal2 s 8442 25225 8550 25335 4 gnd
port 517 nsew
rlabel metal2 s 13914 199 14022 275 4 gnd
port 517 nsew
rlabel metal2 s 18426 21055 18534 21131 4 gnd
port 517 nsew
rlabel metal2 s 5178 1779 5286 1855 4 gnd
port 517 nsew
rlabel metal2 s 15930 7055 16038 7165 4 gnd
port 517 nsew
rlabel metal2 s 8442 12839 8550 12915 4 gnd
port 517 nsew
rlabel metal2 s 8442 12585 8550 12695 4 gnd
port 517 nsew
rlabel metal2 s 8442 19475 8550 19551 4 gnd
port 517 nsew
rlabel metal2 s 8442 10469 8550 10545 4 gnd
port 517 nsew
rlabel metal2 s 15162 21055 15270 21131 4 gnd
port 517 nsew
rlabel metal2 s 7194 515 7302 591 4 gnd
port 517 nsew
rlabel metal2 s 10938 23645 11046 23755 4 gnd
port 517 nsew
rlabel metal2 s 4698 23899 4806 23975 4 gnd
port 517 nsew
rlabel metal2 s 2682 12049 2790 12125 4 gnd
port 517 nsew
rlabel metal2 s 5178 8889 5286 8965 4 gnd
port 517 nsew
rlabel metal2 s 8442 14955 8550 15065 4 gnd
port 517 nsew
rlabel metal2 s 15162 18369 15270 18445 4 gnd
port 517 nsew
rlabel metal2 s 2682 10785 2790 10861 4 gnd
port 517 nsew
rlabel metal2 s 3450 10469 3558 10545 4 gnd
port 517 nsew
rlabel metal2 s 7674 17325 7782 17435 4 gnd
port 517 nsew
rlabel metal2 s 16410 22065 16518 22175 4 gnd
port 517 nsew
rlabel metal2 s 17178 18369 17286 18445 4 gnd
port 517 nsew
rlabel metal2 s 19674 12365 19782 12441 4 gnd
port 517 nsew
rlabel metal2 s 1434 2885 1542 2961 4 gnd
port 517 nsew
rlabel metal2 s 7194 24689 7302 24765 4 gnd
port 517 nsew
rlabel metal2 s 13914 6045 14022 6121 4 gnd
port 517 nsew
rlabel metal2 s 18426 15745 18534 15855 4 gnd
port 517 nsew
rlabel metal2 s 15162 13375 15270 13485 4 gnd
port 517 nsew
rlabel metal2 s 15162 25005 15270 25081 4 gnd
port 517 nsew
rlabel metal2 s 17658 5475 17766 5585 4 gnd
port 517 nsew
rlabel metal2 s 3450 6045 3558 6121 4 gnd
port 517 nsew
rlabel metal2 s 3930 15525 4038 15601 4 gnd
port 517 nsew
rlabel metal2 s 2682 13155 2790 13231 4 gnd
port 517 nsew
rlabel metal2 s 17658 25005 17766 25081 4 gnd
port 517 nsew
rlabel metal2 s 5946 20265 6054 20341 4 gnd
port 517 nsew
rlabel metal2 s 186 7055 294 7165 4 gnd
port 517 nsew
rlabel metal2 s 10170 7845 10278 7955 4 gnd
port 517 nsew
rlabel metal2 s 13434 6519 13542 6595 4 gnd
port 517 nsew
rlabel metal2 s 17658 8415 17766 8491 4 gnd
port 517 nsew
rlabel metal2 s 18426 17895 18534 17971 4 gnd
port 517 nsew
rlabel metal2 s 12666 14419 12774 14495 4 gnd
port 517 nsew
rlabel metal2 s 3930 19949 4038 20025 4 gnd
port 517 nsew
rlabel metal2 s 3450 21845 3558 21921 4 gnd
port 517 nsew
rlabel metal2 s 9690 21055 9798 21131 4 gnd
port 517 nsew
rlabel metal2 s 19674 15999 19782 16075 4 gnd
port 517 nsew
rlabel metal2 s 4698 1305 4806 1381 4 gnd
port 517 nsew
rlabel metal2 s 12666 7845 12774 7955 4 gnd
port 517 nsew
rlabel metal2 s 18426 6519 18534 6595 4 gnd
port 517 nsew
rlabel metal2 s 1434 -55 1542 55 4 gnd
port 517 nsew
rlabel metal2 s 18906 25225 19014 25335 4 gnd
port 517 nsew
rlabel metal2 s 19674 13945 19782 14021 4 gnd
port 517 nsew
rlabel metal2 s 8442 7055 8550 7165 4 gnd
port 517 nsew
rlabel metal2 s 1434 17325 1542 17435 4 gnd
port 517 nsew
rlabel metal2 s 11418 2569 11526 2645 4 gnd
port 517 nsew
rlabel metal2 s 18426 6835 18534 6911 4 gnd
port 517 nsew
rlabel metal2 s 14682 5475 14790 5585 4 gnd
port 517 nsew
rlabel metal2 s 18906 3675 19014 3751 4 gnd
port 517 nsew
rlabel metal2 s 7674 19949 7782 20025 4 gnd
port 517 nsew
rlabel metal2 s 16410 23109 16518 23185 4 gnd
port 517 nsew
rlabel metal2 s 11418 19695 11526 19805 4 gnd
port 517 nsew
rlabel metal2 s 18426 9205 18534 9281 4 gnd
port 517 nsew
rlabel metal2 s 13914 22319 14022 22395 4 gnd
port 517 nsew
rlabel metal2 s 2202 19475 2310 19551 4 gnd
port 517 nsew
rlabel metal2 s 7674 24435 7782 24545 4 gnd
port 517 nsew
rlabel metal2 s 5178 19949 5286 20025 4 gnd
port 517 nsew
rlabel metal2 s 8922 4939 9030 5015 4 gnd
port 517 nsew
rlabel metal2 s 1434 7845 1542 7955 4 gnd
port 517 nsew
rlabel metal2 s 13434 7309 13542 7385 4 gnd
port 517 nsew
rlabel metal2 s 19674 2885 19782 2961 4 gnd
port 517 nsew
rlabel metal2 s 3450 5255 3558 5331 4 gnd
port 517 nsew
rlabel metal2 s 13434 1779 13542 1855 4 gnd
port 517 nsew
rlabel metal2 s 15930 13375 16038 13485 4 gnd
port 517 nsew
rlabel metal2 s 2202 735 2310 845 4 gnd
port 517 nsew
rlabel metal2 s 186 11575 294 11651 4 gnd
port 517 nsew
rlabel metal2 s 5178 15525 5286 15601 4 gnd
port 517 nsew
rlabel metal2 s 4698 18685 4806 18761 4 gnd
port 517 nsew
rlabel metal2 s 8922 11259 9030 11335 4 gnd
port 517 nsew
rlabel metal2 s 17658 -55 17766 55 4 gnd
port 517 nsew
rlabel metal2 s 14682 22855 14790 22965 4 gnd
port 517 nsew
rlabel metal2 s 9690 22319 9798 22395 4 gnd
port 517 nsew
rlabel metal2 s 15162 22319 15270 22395 4 gnd
port 517 nsew
rlabel metal2 s 17658 22855 17766 22965 4 gnd
port 517 nsew
rlabel metal2 s 8442 7845 8550 7955 4 gnd
port 517 nsew
rlabel metal2 s 14682 24435 14790 24545 4 gnd
port 517 nsew
rlabel metal2 s 10938 12585 11046 12695 4 gnd
port 517 nsew
rlabel metal2 s 5946 4149 6054 4225 4 gnd
port 517 nsew
rlabel metal2 s 15930 7845 16038 7955 4 gnd
port 517 nsew
rlabel metal2 s 3930 2315 4038 2425 4 gnd
port 517 nsew
rlabel metal2 s 15930 19159 16038 19235 4 gnd
port 517 nsew
rlabel metal2 s 13434 8889 13542 8965 4 gnd
port 517 nsew
rlabel metal2 s 15930 19949 16038 20025 4 gnd
port 517 nsew
rlabel metal2 s 15930 3359 16038 3435 4 gnd
port 517 nsew
rlabel metal2 s 15162 9995 15270 10071 4 gnd
port 517 nsew
rlabel metal2 s 954 16789 1062 16865 4 gnd
port 517 nsew
rlabel metal2 s 9690 23645 9798 23755 4 gnd
port 517 nsew
rlabel metal2 s 17178 17895 17286 17971 4 gnd
port 517 nsew
rlabel metal2 s 15162 10785 15270 10861 4 gnd
port 517 nsew
rlabel metal2 s 6426 12839 6534 12915 4 gnd
port 517 nsew
rlabel metal2 s 13914 15209 14022 15285 4 gnd
port 517 nsew
rlabel metal2 s 19674 4465 19782 4541 4 gnd
port 517 nsew
rlabel metal2 s 18906 13375 19014 13485 4 gnd
port 517 nsew
rlabel metal2 s 186 22319 294 22395 4 gnd
port 517 nsew
rlabel metal2 s 18906 19949 19014 20025 4 gnd
port 517 nsew
rlabel metal2 s 11418 9995 11526 10071 4 gnd
port 517 nsew
rlabel metal2 s 3450 735 3558 845 4 gnd
port 517 nsew
rlabel metal2 s 8442 23109 8550 23185 4 gnd
port 517 nsew
rlabel metal2 s 18906 22319 19014 22395 4 gnd
port 517 nsew
rlabel metal2 s 15162 11259 15270 11335 4 gnd
port 517 nsew
rlabel metal2 s 11418 16535 11526 16645 4 gnd
port 517 nsew
rlabel metal2 s 5178 9995 5286 10071 4 gnd
port 517 nsew
rlabel metal2 s 10938 4939 11046 5015 4 gnd
port 517 nsew
rlabel metal2 s 16410 5475 16518 5585 4 gnd
port 517 nsew
rlabel metal2 s 12666 3359 12774 3435 4 gnd
port 517 nsew
rlabel metal2 s 13434 8635 13542 8745 4 gnd
port 517 nsew
rlabel metal2 s 186 13629 294 13705 4 gnd
port 517 nsew
rlabel metal2 s 954 24689 1062 24765 4 gnd
port 517 nsew
rlabel metal2 s 18426 21845 18534 21921 4 gnd
port 517 nsew
rlabel metal2 s 19674 24215 19782 24291 4 gnd
port 517 nsew
rlabel metal2 s 1434 23899 1542 23975 4 gnd
port 517 nsew
rlabel metal2 s 5178 21845 5286 21921 4 gnd
port 517 nsew
rlabel metal2 s 13434 11575 13542 11651 4 gnd
port 517 nsew
rlabel metal2 s 13914 9995 14022 10071 4 gnd
port 517 nsew
rlabel metal2 s 15162 10469 15270 10545 4 gnd
port 517 nsew
rlabel metal2 s 11418 1525 11526 1635 4 gnd
port 517 nsew
rlabel metal2 s 13914 14419 14022 14495 4 gnd
port 517 nsew
rlabel metal2 s 15930 11259 16038 11335 4 gnd
port 517 nsew
rlabel metal2 s 13914 21845 14022 21921 4 gnd
port 517 nsew
rlabel metal2 s 3930 5475 4038 5585 4 gnd
port 517 nsew
rlabel metal2 s 18906 23425 19014 23501 4 gnd
port 517 nsew
rlabel metal2 s 8922 18369 9030 18445 4 gnd
port 517 nsew
rlabel metal2 s 15162 14419 15270 14495 4 gnd
port 517 nsew
rlabel metal2 s 18906 10215 19014 10325 4 gnd
port 517 nsew
rlabel metal2 s 13434 7625 13542 7701 4 gnd
port 517 nsew
rlabel metal2 s 7674 7625 7782 7701 4 gnd
port 517 nsew
rlabel metal2 s 13914 22065 14022 22175 4 gnd
port 517 nsew
rlabel metal2 s 7194 1305 7302 1381 4 gnd
port 517 nsew
rlabel metal2 s 5178 3105 5286 3215 4 gnd
port 517 nsew
rlabel metal2 s 8922 14165 9030 14275 4 gnd
port 517 nsew
rlabel metal2 s 12666 6045 12774 6121 4 gnd
port 517 nsew
rlabel metal2 s 4698 5475 4806 5585 4 gnd
port 517 nsew
rlabel metal2 s 10170 14419 10278 14495 4 gnd
port 517 nsew
rlabel metal2 s 4698 22065 4806 22175 4 gnd
port 517 nsew
rlabel metal2 s 16410 16789 16518 16865 4 gnd
port 517 nsew
rlabel metal2 s 8922 19475 9030 19551 4 gnd
port 517 nsew
rlabel metal2 s 18426 15525 18534 15601 4 gnd
port 517 nsew
rlabel metal2 s 6426 10215 6534 10325 4 gnd
port 517 nsew
rlabel metal2 s 186 12049 294 12125 4 gnd
port 517 nsew
rlabel metal2 s 5946 735 6054 845 4 gnd
port 517 nsew
rlabel metal2 s 12186 18369 12294 18445 4 gnd
port 517 nsew
rlabel metal2 s 15162 7055 15270 7165 4 gnd
port 517 nsew
rlabel metal2 s 13434 15209 13542 15285 4 gnd
port 517 nsew
rlabel metal2 s 3930 6045 4038 6121 4 gnd
port 517 nsew
rlabel metal2 s 9690 9205 9798 9281 4 gnd
port 517 nsew
rlabel metal2 s 15162 5475 15270 5585 4 gnd
port 517 nsew
rlabel metal2 s 18426 2885 18534 2961 4 gnd
port 517 nsew
rlabel metal2 s 14682 23109 14790 23185 4 gnd
port 517 nsew
rlabel metal2 s 954 17895 1062 17971 4 gnd
port 517 nsew
rlabel metal2 s 2682 5255 2790 5331 4 gnd
port 517 nsew
rlabel metal2 s 954 1305 1062 1381 4 gnd
port 517 nsew
rlabel metal2 s 2202 20265 2310 20341 4 gnd
port 517 nsew
rlabel metal2 s 17658 23109 17766 23185 4 gnd
port 517 nsew
rlabel metal2 s 4698 10469 4806 10545 4 gnd
port 517 nsew
rlabel metal2 s 7674 18115 7782 18225 4 gnd
port 517 nsew
rlabel metal2 s 6426 19695 6534 19805 4 gnd
port 517 nsew
rlabel metal2 s 3450 7845 3558 7955 4 gnd
port 517 nsew
rlabel metal2 s 2682 5475 2790 5585 4 gnd
port 517 nsew
rlabel metal2 s 7194 23425 7302 23501 4 gnd
port 517 nsew
rlabel metal2 s 13914 8415 14022 8491 4 gnd
port 517 nsew
rlabel metal2 s 6426 21529 6534 21605 4 gnd
port 517 nsew
rlabel metal2 s 10170 735 10278 845 4 gnd
port 517 nsew
rlabel metal2 s 6426 20265 6534 20341 4 gnd
port 517 nsew
rlabel metal2 s 1434 12049 1542 12125 4 gnd
port 517 nsew
rlabel metal2 s 10170 17895 10278 17971 4 gnd
port 517 nsew
rlabel metal2 s 3930 23899 4038 23975 4 gnd
port 517 nsew
rlabel metal2 s 12666 14955 12774 15065 4 gnd
port 517 nsew
rlabel metal2 s 5178 17579 5286 17655 4 gnd
port 517 nsew
rlabel metal2 s 17178 23109 17286 23185 4 gnd
port 517 nsew
rlabel metal2 s 5946 23109 6054 23185 4 gnd
port 517 nsew
rlabel metal2 s 19674 9205 19782 9281 4 gnd
port 517 nsew
rlabel metal2 s 7674 5255 7782 5331 4 gnd
port 517 nsew
rlabel metal2 s 8922 6045 9030 6121 4 gnd
port 517 nsew
rlabel metal2 s 17178 6519 17286 6595 4 gnd
port 517 nsew
rlabel metal2 s 12666 21055 12774 21131 4 gnd
port 517 nsew
rlabel metal2 s 14682 11005 14790 11115 4 gnd
port 517 nsew
rlabel metal2 s 18906 8889 19014 8965 4 gnd
port 517 nsew
rlabel metal2 s 6426 22065 6534 22175 4 gnd
port 517 nsew
rlabel metal2 s 9690 13375 9798 13485 4 gnd
port 517 nsew
rlabel metal2 s 3450 23425 3558 23501 4 gnd
port 517 nsew
rlabel metal2 s 19674 13629 19782 13705 4 gnd
port 517 nsew
rlabel metal2 s 17178 11005 17286 11115 4 gnd
port 517 nsew
rlabel metal2 s 186 24435 294 24545 4 gnd
port 517 nsew
rlabel metal2 s 7194 22065 7302 22175 4 gnd
port 517 nsew
rlabel metal2 s 18906 989 19014 1065 4 gnd
port 517 nsew
rlabel metal2 s 3930 8635 4038 8745 4 gnd
port 517 nsew
rlabel metal2 s 5178 10215 5286 10325 4 gnd
port 517 nsew
rlabel metal2 s 16410 12585 16518 12695 4 gnd
port 517 nsew
rlabel metal2 s 19674 14165 19782 14275 4 gnd
port 517 nsew
rlabel metal2 s 8442 1525 8550 1635 4 gnd
port 517 nsew
rlabel metal2 s 3930 18905 4038 19015 4 gnd
port 517 nsew
rlabel metal2 s 8442 13375 8550 13485 4 gnd
port 517 nsew
rlabel metal2 s 1434 11795 1542 11905 4 gnd
port 517 nsew
rlabel metal2 s 3450 18905 3558 19015 4 gnd
port 517 nsew
rlabel metal2 s 10170 11005 10278 11115 4 gnd
port 517 nsew
rlabel metal2 s 19674 10469 19782 10545 4 gnd
port 517 nsew
rlabel metal2 s 15930 21529 16038 21605 4 gnd
port 517 nsew
rlabel metal2 s 7194 13629 7302 13705 4 gnd
port 517 nsew
rlabel metal2 s 7194 1779 7302 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 8415 7782 8491 4 gnd
port 517 nsew
rlabel metal2 s 18426 5729 18534 5805 4 gnd
port 517 nsew
rlabel metal2 s 8922 20265 9030 20341 4 gnd
port 517 nsew
rlabel metal2 s 954 2885 1062 2961 4 gnd
port 517 nsew
rlabel metal2 s 4698 21275 4806 21385 4 gnd
port 517 nsew
rlabel metal2 s 8922 16535 9030 16645 4 gnd
port 517 nsew
rlabel metal2 s 10938 23425 11046 23501 4 gnd
port 517 nsew
rlabel metal2 s 13914 8635 14022 8745 4 gnd
port 517 nsew
rlabel metal2 s 14682 12585 14790 12695 4 gnd
port 517 nsew
rlabel metal2 s 17178 5475 17286 5585 4 gnd
port 517 nsew
rlabel metal2 s 3930 24215 4038 24291 4 gnd
port 517 nsew
rlabel metal2 s 8922 735 9030 845 4 gnd
port 517 nsew
rlabel metal2 s 954 13155 1062 13231 4 gnd
port 517 nsew
rlabel metal2 s 16410 -55 16518 55 4 gnd
port 517 nsew
rlabel metal2 s 12666 16789 12774 16865 4 gnd
port 517 nsew
rlabel metal2 s 1434 20265 1542 20341 4 gnd
port 517 nsew
rlabel metal2 s 15162 16789 15270 16865 4 gnd
port 517 nsew
rlabel metal2 s 14682 7055 14790 7165 4 gnd
port 517 nsew
rlabel metal2 s 5178 14955 5286 15065 4 gnd
port 517 nsew
rlabel metal2 s 3450 9205 3558 9281 4 gnd
port 517 nsew
rlabel metal2 s 8442 21055 8550 21131 4 gnd
port 517 nsew
rlabel metal2 s 18426 22065 18534 22175 4 gnd
port 517 nsew
rlabel metal2 s 13434 21845 13542 21921 4 gnd
port 517 nsew
rlabel metal2 s 2202 9679 2310 9755 4 gnd
port 517 nsew
rlabel metal2 s 2682 7055 2790 7165 4 gnd
port 517 nsew
rlabel metal2 s 3450 17105 3558 17181 4 gnd
port 517 nsew
rlabel metal2 s 7674 15999 7782 16075 4 gnd
port 517 nsew
rlabel metal2 s 7194 24215 7302 24291 4 gnd
port 517 nsew
rlabel metal2 s 18426 735 18534 845 4 gnd
port 517 nsew
rlabel metal2 s 2202 8099 2310 8175 4 gnd
port 517 nsew
rlabel metal2 s 4698 1525 4806 1635 4 gnd
port 517 nsew
rlabel metal2 s 9690 3105 9798 3215 4 gnd
port 517 nsew
rlabel metal2 s 13434 16315 13542 16391 4 gnd
port 517 nsew
rlabel metal2 s 6426 13629 6534 13705 4 gnd
port 517 nsew
rlabel metal2 s 8442 1779 8550 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 18369 7782 18445 4 gnd
port 517 nsew
rlabel metal2 s 14682 14955 14790 15065 4 gnd
port 517 nsew
rlabel metal2 s 13914 25005 14022 25081 4 gnd
port 517 nsew
rlabel metal2 s 1434 12365 1542 12441 4 gnd
port 517 nsew
rlabel metal2 s 6426 23899 6534 23975 4 gnd
port 517 nsew
rlabel metal2 s 4698 17105 4806 17181 4 gnd
port 517 nsew
rlabel metal2 s 5946 16535 6054 16645 4 gnd
port 517 nsew
rlabel metal2 s 3450 12365 3558 12441 4 gnd
port 517 nsew
rlabel metal2 s 8922 19949 9030 20025 4 gnd
port 517 nsew
rlabel metal2 s 13434 21275 13542 21385 4 gnd
port 517 nsew
rlabel metal2 s 8922 24689 9030 24765 4 gnd
port 517 nsew
rlabel metal2 s 17658 15745 17766 15855 4 gnd
port 517 nsew
rlabel metal2 s 1434 17579 1542 17655 4 gnd
port 517 nsew
rlabel metal2 s 19674 21275 19782 21385 4 gnd
port 517 nsew
rlabel metal2 s 11418 12585 11526 12695 4 gnd
port 517 nsew
rlabel metal2 s 13434 12049 13542 12125 4 gnd
port 517 nsew
rlabel metal2 s 3450 6835 3558 6911 4 gnd
port 517 nsew
rlabel metal2 s 13434 21529 13542 21605 4 gnd
port 517 nsew
rlabel metal2 s 15930 5255 16038 5331 4 gnd
port 517 nsew
rlabel metal2 s 16410 19475 16518 19551 4 gnd
port 517 nsew
rlabel metal2 s 17658 11259 17766 11335 4 gnd
port 517 nsew
rlabel metal2 s 18906 8099 19014 8175 4 gnd
port 517 nsew
rlabel metal2 s 14682 25005 14790 25081 4 gnd
port 517 nsew
rlabel metal2 s 19674 14955 19782 15065 4 gnd
port 517 nsew
rlabel metal2 s 6426 8889 6534 8965 4 gnd
port 517 nsew
rlabel metal2 s 2202 16315 2310 16391 4 gnd
port 517 nsew
rlabel metal2 s 16410 17579 16518 17655 4 gnd
port 517 nsew
rlabel metal2 s 19674 20485 19782 20595 4 gnd
port 517 nsew
rlabel metal2 s 17178 23645 17286 23755 4 gnd
port 517 nsew
rlabel metal2 s 3930 12839 4038 12915 4 gnd
port 517 nsew
rlabel metal2 s 8922 3105 9030 3215 4 gnd
port 517 nsew
rlabel metal2 s 12186 19695 12294 19805 4 gnd
port 517 nsew
rlabel metal2 s 8922 16315 9030 16391 4 gnd
port 517 nsew
rlabel metal2 s 8922 22065 9030 22175 4 gnd
port 517 nsew
rlabel metal2 s 5178 21529 5286 21605 4 gnd
port 517 nsew
rlabel metal2 s 7674 515 7782 591 4 gnd
port 517 nsew
rlabel metal2 s 4698 14419 4806 14495 4 gnd
port 517 nsew
rlabel metal2 s 3450 22855 3558 22965 4 gnd
port 517 nsew
rlabel metal2 s 17658 21055 17766 21131 4 gnd
port 517 nsew
rlabel metal2 s 8922 21275 9030 21385 4 gnd
port 517 nsew
rlabel metal2 s 10170 15209 10278 15285 4 gnd
port 517 nsew
rlabel metal2 s 15930 6835 16038 6911 4 gnd
port 517 nsew
rlabel metal2 s 15162 11795 15270 11905 4 gnd
port 517 nsew
rlabel metal2 s 8442 18905 8550 19015 4 gnd
port 517 nsew
rlabel metal2 s 4698 22635 4806 22711 4 gnd
port 517 nsew
rlabel metal2 s 6426 25005 6534 25081 4 gnd
port 517 nsew
rlabel metal2 s 1434 15999 1542 16075 4 gnd
port 517 nsew
rlabel metal2 s 9690 9679 9798 9755 4 gnd
port 517 nsew
rlabel metal2 s 17658 24215 17766 24291 4 gnd
port 517 nsew
rlabel metal2 s 9690 25005 9798 25081 4 gnd
port 517 nsew
rlabel metal2 s 2202 9995 2310 10071 4 gnd
port 517 nsew
rlabel metal2 s 954 8099 1062 8175 4 gnd
port 517 nsew
rlabel metal2 s 12186 18685 12294 18761 4 gnd
port 517 nsew
rlabel metal2 s 8922 22635 9030 22711 4 gnd
port 517 nsew
rlabel metal2 s 15162 21529 15270 21605 4 gnd
port 517 nsew
rlabel metal2 s 954 11795 1062 11905 4 gnd
port 517 nsew
rlabel metal2 s 8442 7309 8550 7385 4 gnd
port 517 nsew
rlabel metal2 s 8442 19949 8550 20025 4 gnd
port 517 nsew
rlabel metal2 s 16410 4149 16518 4225 4 gnd
port 517 nsew
rlabel metal2 s 5946 15745 6054 15855 4 gnd
port 517 nsew
rlabel metal2 s 10938 12365 11046 12441 4 gnd
port 517 nsew
rlabel metal2 s 2682 6265 2790 6375 4 gnd
port 517 nsew
rlabel metal2 s 10938 13945 11046 14021 4 gnd
port 517 nsew
rlabel metal2 s 12186 22855 12294 22965 4 gnd
port 517 nsew
rlabel metal2 s 14682 735 14790 845 4 gnd
port 517 nsew
rlabel metal2 s 18426 14955 18534 15065 4 gnd
port 517 nsew
rlabel metal2 s 5178 16535 5286 16645 4 gnd
port 517 nsew
rlabel metal2 s 17178 7309 17286 7385 4 gnd
port 517 nsew
rlabel metal2 s 12666 21529 12774 21605 4 gnd
port 517 nsew
rlabel metal2 s 7194 9679 7302 9755 4 gnd
port 517 nsew
rlabel metal2 s 9690 24435 9798 24545 4 gnd
port 517 nsew
rlabel metal2 s 186 17895 294 17971 4 gnd
port 517 nsew
rlabel metal2 s 186 3895 294 4005 4 gnd
port 517 nsew
rlabel metal2 s 12186 8415 12294 8491 4 gnd
port 517 nsew
rlabel metal2 s 18906 -55 19014 55 4 gnd
port 517 nsew
rlabel metal2 s 19674 21529 19782 21605 4 gnd
port 517 nsew
rlabel metal2 s 18906 4939 19014 5015 4 gnd
port 517 nsew
rlabel metal2 s 2202 13945 2310 14021 4 gnd
port 517 nsew
rlabel metal2 s 2682 3105 2790 3215 4 gnd
port 517 nsew
rlabel metal2 s 11418 6519 11526 6595 4 gnd
port 517 nsew
rlabel metal2 s 10938 989 11046 1065 4 gnd
port 517 nsew
rlabel metal2 s 7194 13945 7302 14021 4 gnd
port 517 nsew
rlabel metal2 s 4698 15999 4806 16075 4 gnd
port 517 nsew
rlabel metal2 s 4698 16789 4806 16865 4 gnd
port 517 nsew
rlabel metal2 s 12666 9679 12774 9755 4 gnd
port 517 nsew
rlabel metal2 s 14682 20739 14790 20815 4 gnd
port 517 nsew
rlabel metal2 s 6426 6045 6534 6121 4 gnd
port 517 nsew
rlabel metal2 s 15162 15525 15270 15601 4 gnd
port 517 nsew
rlabel metal2 s 5178 -55 5286 55 4 gnd
port 517 nsew
rlabel metal2 s 14682 2315 14790 2425 4 gnd
port 517 nsew
rlabel metal2 s 16410 18115 16518 18225 4 gnd
port 517 nsew
rlabel metal2 s 1434 15745 1542 15855 4 gnd
port 517 nsew
rlabel metal2 s 12666 2885 12774 2961 4 gnd
port 517 nsew
rlabel metal2 s 186 15525 294 15601 4 gnd
port 517 nsew
rlabel metal2 s 7194 15209 7302 15285 4 gnd
port 517 nsew
rlabel metal2 s 19674 15209 19782 15285 4 gnd
port 517 nsew
rlabel metal2 s 954 23899 1062 23975 4 gnd
port 517 nsew
rlabel metal2 s 18426 11005 18534 11115 4 gnd
port 517 nsew
rlabel metal2 s 7194 19159 7302 19235 4 gnd
port 517 nsew
rlabel metal2 s 186 4465 294 4541 4 gnd
port 517 nsew
rlabel metal2 s 2682 11259 2790 11335 4 gnd
port 517 nsew
rlabel metal2 s 17178 4465 17286 4541 4 gnd
port 517 nsew
rlabel metal2 s 11418 4685 11526 4795 4 gnd
port 517 nsew
rlabel metal2 s 11418 11795 11526 11905 4 gnd
port 517 nsew
rlabel metal2 s 18906 17105 19014 17181 4 gnd
port 517 nsew
rlabel metal2 s 5178 12365 5286 12441 4 gnd
port 517 nsew
rlabel metal2 s 7674 19475 7782 19551 4 gnd
port 517 nsew
rlabel metal2 s 12186 735 12294 845 4 gnd
port 517 nsew
rlabel metal2 s 17178 24215 17286 24291 4 gnd
port 517 nsew
rlabel metal2 s 18426 20265 18534 20341 4 gnd
port 517 nsew
rlabel metal2 s 19674 11575 19782 11651 4 gnd
port 517 nsew
rlabel metal2 s 6426 8635 6534 8745 4 gnd
port 517 nsew
rlabel metal2 s 8442 19695 8550 19805 4 gnd
port 517 nsew
rlabel metal2 s 5178 7055 5286 7165 4 gnd
port 517 nsew
rlabel metal2 s 19674 21845 19782 21921 4 gnd
port 517 nsew
rlabel metal2 s 186 12839 294 12915 4 gnd
port 517 nsew
rlabel metal2 s 16410 18905 16518 19015 4 gnd
port 517 nsew
rlabel metal2 s 17178 19949 17286 20025 4 gnd
port 517 nsew
rlabel metal2 s 3930 22065 4038 22175 4 gnd
port 517 nsew
rlabel metal2 s 3450 22065 3558 22175 4 gnd
port 517 nsew
rlabel metal2 s 17658 2569 17766 2645 4 gnd
port 517 nsew
rlabel metal2 s 15162 13945 15270 14021 4 gnd
port 517 nsew
rlabel metal2 s 186 8415 294 8491 4 gnd
port 517 nsew
rlabel metal2 s 2202 15999 2310 16075 4 gnd
port 517 nsew
rlabel metal2 s 12186 3675 12294 3751 4 gnd
port 517 nsew
rlabel metal2 s 14682 3105 14790 3215 4 gnd
port 517 nsew
rlabel metal2 s 3450 4465 3558 4541 4 gnd
port 517 nsew
rlabel metal2 s 17658 18369 17766 18445 4 gnd
port 517 nsew
rlabel metal2 s 3930 19475 4038 19551 4 gnd
port 517 nsew
rlabel metal2 s 9690 18115 9798 18225 4 gnd
port 517 nsew
rlabel metal2 s 2202 10215 2310 10325 4 gnd
port 517 nsew
rlabel metal2 s 17178 9205 17286 9281 4 gnd
port 517 nsew
rlabel metal2 s 15162 8635 15270 8745 4 gnd
port 517 nsew
rlabel metal2 s 18906 11005 19014 11115 4 gnd
port 517 nsew
rlabel metal2 s 15162 7309 15270 7385 4 gnd
port 517 nsew
rlabel metal2 s 5946 2885 6054 2961 4 gnd
port 517 nsew
rlabel metal2 s 1434 13155 1542 13231 4 gnd
port 517 nsew
rlabel metal2 s 13914 21275 14022 21385 4 gnd
port 517 nsew
rlabel metal2 s 7674 21845 7782 21921 4 gnd
port 517 nsew
rlabel metal2 s 954 18369 1062 18445 4 gnd
port 517 nsew
rlabel metal2 s 7674 15525 7782 15601 4 gnd
port 517 nsew
rlabel metal2 s 17178 21529 17286 21605 4 gnd
port 517 nsew
rlabel metal2 s 10170 5475 10278 5585 4 gnd
port 517 nsew
rlabel metal2 s 15162 4465 15270 4541 4 gnd
port 517 nsew
rlabel metal2 s 16410 2315 16518 2425 4 gnd
port 517 nsew
rlabel metal2 s 12666 5729 12774 5805 4 gnd
port 517 nsew
rlabel metal2 s 19674 11259 19782 11335 4 gnd
port 517 nsew
rlabel metal2 s 7674 4685 7782 4795 4 gnd
port 517 nsew
rlabel metal2 s 13914 10469 14022 10545 4 gnd
port 517 nsew
rlabel metal2 s 4698 13629 4806 13705 4 gnd
port 517 nsew
rlabel metal2 s 186 1779 294 1855 4 gnd
port 517 nsew
rlabel metal2 s 16410 5729 16518 5805 4 gnd
port 517 nsew
rlabel metal2 s 5178 18115 5286 18225 4 gnd
port 517 nsew
rlabel metal2 s 5946 19949 6054 20025 4 gnd
port 517 nsew
rlabel metal2 s 17658 17895 17766 17971 4 gnd
port 517 nsew
rlabel metal2 s 1434 10469 1542 10545 4 gnd
port 517 nsew
rlabel metal2 s 2202 17579 2310 17655 4 gnd
port 517 nsew
rlabel metal2 s 17178 4149 17286 4225 4 gnd
port 517 nsew
rlabel metal2 s 10170 12585 10278 12695 4 gnd
port 517 nsew
rlabel metal2 s 186 12585 294 12695 4 gnd
port 517 nsew
rlabel metal2 s 6426 10785 6534 10861 4 gnd
port 517 nsew
rlabel metal2 s 3930 11575 4038 11651 4 gnd
port 517 nsew
rlabel metal2 s 4698 6835 4806 6911 4 gnd
port 517 nsew
rlabel metal2 s 18426 11575 18534 11651 4 gnd
port 517 nsew
rlabel metal2 s 13434 21055 13542 21131 4 gnd
port 517 nsew
rlabel metal2 s 18426 11259 18534 11335 4 gnd
port 517 nsew
rlabel metal2 s 13434 4939 13542 5015 4 gnd
port 517 nsew
rlabel metal2 s 13914 3359 14022 3435 4 gnd
port 517 nsew
rlabel metal2 s 5178 2315 5286 2425 4 gnd
port 517 nsew
rlabel metal2 s 17658 20265 17766 20341 4 gnd
port 517 nsew
rlabel metal2 s 17178 7845 17286 7955 4 gnd
port 517 nsew
rlabel metal2 s 8442 10785 8550 10861 4 gnd
port 517 nsew
rlabel metal2 s 4698 20485 4806 20595 4 gnd
port 517 nsew
rlabel metal2 s 2682 4465 2790 4541 4 gnd
port 517 nsew
rlabel metal2 s 5178 22065 5286 22175 4 gnd
port 517 nsew
rlabel metal2 s 8922 25005 9030 25081 4 gnd
port 517 nsew
rlabel metal2 s 10170 5255 10278 5331 4 gnd
port 517 nsew
rlabel metal2 s 7194 3675 7302 3751 4 gnd
port 517 nsew
rlabel metal2 s 10938 16535 11046 16645 4 gnd
port 517 nsew
rlabel metal2 s 13914 13629 14022 13705 4 gnd
port 517 nsew
rlabel metal2 s 14682 17325 14790 17435 4 gnd
port 517 nsew
rlabel metal2 s 6426 3895 6534 4005 4 gnd
port 517 nsew
rlabel metal2 s 7674 7309 7782 7385 4 gnd
port 517 nsew
rlabel metal2 s 2682 16789 2790 16865 4 gnd
port 517 nsew
rlabel metal2 s 10170 18115 10278 18225 4 gnd
port 517 nsew
rlabel metal2 s 12666 989 12774 1065 4 gnd
port 517 nsew
rlabel metal2 s 18906 18115 19014 18225 4 gnd
port 517 nsew
rlabel metal2 s 10938 2095 11046 2171 4 gnd
port 517 nsew
rlabel metal2 s 15930 1305 16038 1381 4 gnd
port 517 nsew
rlabel metal2 s 15162 15745 15270 15855 4 gnd
port 517 nsew
rlabel metal2 s 1434 18369 1542 18445 4 gnd
port 517 nsew
rlabel metal2 s 13914 735 14022 845 4 gnd
port 517 nsew
rlabel metal2 s 2202 3359 2310 3435 4 gnd
port 517 nsew
rlabel metal2 s 19674 3359 19782 3435 4 gnd
port 517 nsew
rlabel metal2 s 14682 1305 14790 1381 4 gnd
port 517 nsew
rlabel metal2 s 7194 9995 7302 10071 4 gnd
port 517 nsew
rlabel metal2 s 17658 515 17766 591 4 gnd
port 517 nsew
rlabel metal2 s 7194 4149 7302 4225 4 gnd
port 517 nsew
rlabel metal2 s 1434 23109 1542 23185 4 gnd
port 517 nsew
rlabel metal2 s 13914 8099 14022 8175 4 gnd
port 517 nsew
rlabel metal2 s 15162 23109 15270 23185 4 gnd
port 517 nsew
rlabel metal2 s 8442 15209 8550 15285 4 gnd
port 517 nsew
rlabel metal2 s 1434 6045 1542 6121 4 gnd
port 517 nsew
rlabel metal2 s 8442 22065 8550 22175 4 gnd
port 517 nsew
rlabel metal2 s 14682 9679 14790 9755 4 gnd
port 517 nsew
rlabel metal2 s 17178 20739 17286 20815 4 gnd
port 517 nsew
rlabel metal2 s 3450 1779 3558 1855 4 gnd
port 517 nsew
rlabel metal2 s 3930 18685 4038 18761 4 gnd
port 517 nsew
rlabel metal2 s 8922 8415 9030 8491 4 gnd
port 517 nsew
rlabel metal2 s 3450 23899 3558 23975 4 gnd
port 517 nsew
rlabel metal2 s 5946 13375 6054 13485 4 gnd
port 517 nsew
rlabel metal2 s 11418 19949 11526 20025 4 gnd
port 517 nsew
rlabel metal2 s 7674 10469 7782 10545 4 gnd
port 517 nsew
rlabel metal2 s 954 3675 1062 3751 4 gnd
port 517 nsew
rlabel metal2 s 2202 19159 2310 19235 4 gnd
port 517 nsew
rlabel metal2 s 3930 18369 4038 18445 4 gnd
port 517 nsew
rlabel metal2 s 16410 7055 16518 7165 4 gnd
port 517 nsew
rlabel metal2 s 16410 8635 16518 8745 4 gnd
port 517 nsew
rlabel metal2 s 19674 17579 19782 17655 4 gnd
port 517 nsew
rlabel metal2 s 9690 17579 9798 17655 4 gnd
port 517 nsew
rlabel metal2 s 16410 20265 16518 20341 4 gnd
port 517 nsew
rlabel metal2 s 1434 22855 1542 22965 4 gnd
port 517 nsew
rlabel metal2 s 17178 3895 17286 4005 4 gnd
port 517 nsew
rlabel metal2 s 7194 8099 7302 8175 4 gnd
port 517 nsew
rlabel metal2 s 2682 15745 2790 15855 4 gnd
port 517 nsew
rlabel metal2 s 8442 8099 8550 8175 4 gnd
port 517 nsew
rlabel metal2 s 8442 20739 8550 20815 4 gnd
port 517 nsew
rlabel metal2 s 16410 21845 16518 21921 4 gnd
port 517 nsew
rlabel metal2 s 18906 22855 19014 22965 4 gnd
port 517 nsew
rlabel metal2 s 14682 8635 14790 8745 4 gnd
port 517 nsew
rlabel metal2 s 15162 3359 15270 3435 4 gnd
port 517 nsew
rlabel metal2 s 7194 2095 7302 2171 4 gnd
port 517 nsew
rlabel metal2 s 15930 989 16038 1065 4 gnd
port 517 nsew
rlabel metal2 s 11418 22065 11526 22175 4 gnd
port 517 nsew
rlabel metal2 s 10170 13945 10278 14021 4 gnd
port 517 nsew
rlabel metal2 s 1434 22065 1542 22175 4 gnd
port 517 nsew
rlabel metal2 s 16410 18369 16518 18445 4 gnd
port 517 nsew
rlabel metal2 s 14682 6519 14790 6595 4 gnd
port 517 nsew
rlabel metal2 s 3930 199 4038 275 4 gnd
port 517 nsew
rlabel metal2 s 6426 18369 6534 18445 4 gnd
port 517 nsew
rlabel metal2 s 10170 7055 10278 7165 4 gnd
port 517 nsew
rlabel metal2 s 5946 20739 6054 20815 4 gnd
port 517 nsew
rlabel metal2 s 15162 3105 15270 3215 4 gnd
port 517 nsew
rlabel metal2 s 2202 2315 2310 2425 4 gnd
port 517 nsew
rlabel metal2 s 12186 199 12294 275 4 gnd
port 517 nsew
rlabel metal2 s 954 16315 1062 16391 4 gnd
port 517 nsew
rlabel metal2 s 13914 5475 14022 5585 4 gnd
port 517 nsew
rlabel metal2 s 5178 12049 5286 12125 4 gnd
port 517 nsew
rlabel metal2 s 4698 7309 4806 7385 4 gnd
port 517 nsew
rlabel metal2 s 5178 19159 5286 19235 4 gnd
port 517 nsew
rlabel metal2 s 1434 11259 1542 11335 4 gnd
port 517 nsew
rlabel metal2 s 4698 4939 4806 5015 4 gnd
port 517 nsew
rlabel metal2 s 3930 10785 4038 10861 4 gnd
port 517 nsew
rlabel metal2 s 13434 4149 13542 4225 4 gnd
port 517 nsew
rlabel metal2 s 11418 19159 11526 19235 4 gnd
port 517 nsew
rlabel metal2 s 10170 19695 10278 19805 4 gnd
port 517 nsew
rlabel metal2 s 186 19159 294 19235 4 gnd
port 517 nsew
rlabel metal2 s 14682 9995 14790 10071 4 gnd
port 517 nsew
rlabel metal2 s 3450 17895 3558 17971 4 gnd
port 517 nsew
rlabel metal2 s 5946 11795 6054 11905 4 gnd
port 517 nsew
rlabel metal2 s 4698 5255 4806 5331 4 gnd
port 517 nsew
rlabel metal2 s 11418 18115 11526 18225 4 gnd
port 517 nsew
rlabel metal2 s 12186 12585 12294 12695 4 gnd
port 517 nsew
rlabel metal2 s 3450 19949 3558 20025 4 gnd
port 517 nsew
rlabel metal2 s 7674 18685 7782 18761 4 gnd
port 517 nsew
rlabel metal2 s 18906 1779 19014 1855 4 gnd
port 517 nsew
rlabel metal2 s 4698 4465 4806 4541 4 gnd
port 517 nsew
rlabel metal2 s 15930 8099 16038 8175 4 gnd
port 517 nsew
rlabel metal2 s 15930 8889 16038 8965 4 gnd
port 517 nsew
rlabel metal2 s 2682 23425 2790 23501 4 gnd
port 517 nsew
rlabel metal2 s 3930 7309 4038 7385 4 gnd
port 517 nsew
rlabel metal2 s 8442 25005 8550 25081 4 gnd
port 517 nsew
rlabel metal2 s 6426 14735 6534 14811 4 gnd
port 517 nsew
rlabel metal2 s 18426 9425 18534 9535 4 gnd
port 517 nsew
rlabel metal2 s 7674 9995 7782 10071 4 gnd
port 517 nsew
rlabel metal2 s 17178 11795 17286 11905 4 gnd
port 517 nsew
rlabel metal2 s 12666 4939 12774 5015 4 gnd
port 517 nsew
rlabel metal2 s 14682 8889 14790 8965 4 gnd
port 517 nsew
rlabel metal2 s 13434 11259 13542 11335 4 gnd
port 517 nsew
rlabel metal2 s 19674 14735 19782 14811 4 gnd
port 517 nsew
rlabel metal2 s 13914 22855 14022 22965 4 gnd
port 517 nsew
rlabel metal2 s 4698 23425 4806 23501 4 gnd
port 517 nsew
rlabel metal2 s 15162 6265 15270 6375 4 gnd
port 517 nsew
rlabel metal2 s 1434 6835 1542 6911 4 gnd
port 517 nsew
rlabel metal2 s 1434 6519 1542 6595 4 gnd
port 517 nsew
rlabel metal2 s 19674 3675 19782 3751 4 gnd
port 517 nsew
rlabel metal2 s 5946 22065 6054 22175 4 gnd
port 517 nsew
rlabel metal2 s 3450 8889 3558 8965 4 gnd
port 517 nsew
rlabel metal2 s 1434 13945 1542 14021 4 gnd
port 517 nsew
rlabel metal2 s 4698 16535 4806 16645 4 gnd
port 517 nsew
rlabel metal2 s 186 18685 294 18761 4 gnd
port 517 nsew
rlabel metal2 s 8442 15745 8550 15855 4 gnd
port 517 nsew
rlabel metal2 s 1434 8099 1542 8175 4 gnd
port 517 nsew
rlabel metal2 s 186 15209 294 15285 4 gnd
port 517 nsew
rlabel metal2 s 16410 24435 16518 24545 4 gnd
port 517 nsew
rlabel metal2 s 8442 9995 8550 10071 4 gnd
port 517 nsew
rlabel metal2 s 2202 23425 2310 23501 4 gnd
port 517 nsew
rlabel metal2 s 9690 18905 9798 19015 4 gnd
port 517 nsew
rlabel metal2 s 13434 13629 13542 13705 4 gnd
port 517 nsew
rlabel metal2 s 14682 17579 14790 17655 4 gnd
port 517 nsew
rlabel metal2 s 3930 3359 4038 3435 4 gnd
port 517 nsew
rlabel metal2 s 7674 20739 7782 20815 4 gnd
port 517 nsew
rlabel metal2 s 13434 18115 13542 18225 4 gnd
port 517 nsew
rlabel metal2 s 16410 515 16518 591 4 gnd
port 517 nsew
rlabel metal2 s 186 7625 294 7701 4 gnd
port 517 nsew
rlabel metal2 s 10938 24435 11046 24545 4 gnd
port 517 nsew
rlabel metal2 s 954 4149 1062 4225 4 gnd
port 517 nsew
rlabel metal2 s 5178 17105 5286 17181 4 gnd
port 517 nsew
rlabel metal2 s 17178 12365 17286 12441 4 gnd
port 517 nsew
rlabel metal2 s 2202 22855 2310 22965 4 gnd
port 517 nsew
rlabel metal2 s 13914 18685 14022 18761 4 gnd
port 517 nsew
rlabel metal2 s 19674 24689 19782 24765 4 gnd
port 517 nsew
rlabel metal2 s 10938 22065 11046 22175 4 gnd
port 517 nsew
rlabel metal2 s 5946 17105 6054 17181 4 gnd
port 517 nsew
rlabel metal2 s 18426 10215 18534 10325 4 gnd
port 517 nsew
rlabel metal2 s 15162 6045 15270 6121 4 gnd
port 517 nsew
rlabel metal2 s 5178 5475 5286 5585 4 gnd
port 517 nsew
rlabel metal2 s 6426 5475 6534 5585 4 gnd
port 517 nsew
rlabel metal2 s 186 4939 294 5015 4 gnd
port 517 nsew
rlabel metal2 s 15930 14735 16038 14811 4 gnd
port 517 nsew
rlabel metal2 s 11418 18685 11526 18761 4 gnd
port 517 nsew
rlabel metal2 s 13434 515 13542 591 4 gnd
port 517 nsew
rlabel metal2 s 17658 15999 17766 16075 4 gnd
port 517 nsew
rlabel metal2 s 2202 15525 2310 15601 4 gnd
port 517 nsew
rlabel metal2 s 3930 23109 4038 23185 4 gnd
port 517 nsew
rlabel metal2 s 12186 1305 12294 1381 4 gnd
port 517 nsew
rlabel metal2 s 15162 13155 15270 13231 4 gnd
port 517 nsew
rlabel metal2 s 7194 11005 7302 11115 4 gnd
port 517 nsew
rlabel metal2 s 17178 199 17286 275 4 gnd
port 517 nsew
rlabel metal2 s 2682 2569 2790 2645 4 gnd
port 517 nsew
rlabel metal2 s 5178 16315 5286 16391 4 gnd
port 517 nsew
rlabel metal2 s 13434 18369 13542 18445 4 gnd
port 517 nsew
rlabel metal2 s 15162 9205 15270 9281 4 gnd
port 517 nsew
rlabel metal2 s 10938 18369 11046 18445 4 gnd
port 517 nsew
rlabel metal2 s 17658 3895 17766 4005 4 gnd
port 517 nsew
rlabel metal2 s 15162 1305 15270 1381 4 gnd
port 517 nsew
rlabel metal2 s 4698 4149 4806 4225 4 gnd
port 517 nsew
rlabel metal2 s 4698 5729 4806 5805 4 gnd
port 517 nsew
rlabel metal2 s 7674 24215 7782 24291 4 gnd
port 517 nsew
rlabel metal2 s 12666 21845 12774 21921 4 gnd
port 517 nsew
rlabel metal2 s 2202 9205 2310 9281 4 gnd
port 517 nsew
rlabel metal2 s 954 16535 1062 16645 4 gnd
port 517 nsew
rlabel metal2 s 6426 989 6534 1065 4 gnd
port 517 nsew
rlabel metal2 s 18906 24435 19014 24545 4 gnd
port 517 nsew
rlabel metal2 s 11418 13629 11526 13705 4 gnd
port 517 nsew
rlabel metal2 s 6426 14165 6534 14275 4 gnd
port 517 nsew
rlabel metal2 s 12666 10215 12774 10325 4 gnd
port 517 nsew
rlabel metal2 s 7194 25005 7302 25081 4 gnd
port 517 nsew
rlabel metal2 s 15930 22065 16038 22175 4 gnd
port 517 nsew
rlabel metal2 s 10170 5729 10278 5805 4 gnd
port 517 nsew
rlabel metal2 s 19674 14419 19782 14495 4 gnd
port 517 nsew
rlabel metal2 s 10170 17579 10278 17655 4 gnd
port 517 nsew
rlabel metal2 s 16410 20739 16518 20815 4 gnd
port 517 nsew
rlabel metal2 s 3450 2095 3558 2171 4 gnd
port 517 nsew
rlabel metal2 s 10938 3105 11046 3215 4 gnd
port 517 nsew
rlabel metal2 s 10170 14955 10278 15065 4 gnd
port 517 nsew
rlabel metal2 s 13434 19475 13542 19551 4 gnd
port 517 nsew
rlabel metal2 s 186 6045 294 6121 4 gnd
port 517 nsew
rlabel metal2 s 9690 6519 9798 6595 4 gnd
port 517 nsew
rlabel metal2 s 5946 12585 6054 12695 4 gnd
port 517 nsew
rlabel metal2 s 17658 21529 17766 21605 4 gnd
port 517 nsew
rlabel metal2 s 19674 9425 19782 9535 4 gnd
port 517 nsew
rlabel metal2 s 2202 5255 2310 5331 4 gnd
port 517 nsew
rlabel metal2 s 1434 7055 1542 7165 4 gnd
port 517 nsew
rlabel metal2 s 6426 24215 6534 24291 4 gnd
port 517 nsew
rlabel metal2 s 954 4685 1062 4795 4 gnd
port 517 nsew
rlabel metal2 s 8922 989 9030 1065 4 gnd
port 517 nsew
rlabel metal2 s 19674 10215 19782 10325 4 gnd
port 517 nsew
rlabel metal2 s 186 3359 294 3435 4 gnd
port 517 nsew
rlabel metal2 s 5946 14165 6054 14275 4 gnd
port 517 nsew
rlabel metal2 s 19674 9995 19782 10071 4 gnd
port 517 nsew
rlabel metal2 s 10938 14165 11046 14275 4 gnd
port 517 nsew
rlabel metal2 s 1434 199 1542 275 4 gnd
port 517 nsew
rlabel metal2 s 2202 21055 2310 21131 4 gnd
port 517 nsew
rlabel metal2 s 6426 9205 6534 9281 4 gnd
port 517 nsew
rlabel metal2 s 5946 10215 6054 10325 4 gnd
port 517 nsew
rlabel metal2 s 15930 20739 16038 20815 4 gnd
port 517 nsew
rlabel metal2 s 18906 24689 19014 24765 4 gnd
port 517 nsew
rlabel metal2 s 1434 3895 1542 4005 4 gnd
port 517 nsew
rlabel metal2 s 17658 7625 17766 7701 4 gnd
port 517 nsew
rlabel metal2 s 10170 199 10278 275 4 gnd
port 517 nsew
rlabel metal2 s 12186 18905 12294 19015 4 gnd
port 517 nsew
rlabel metal2 s 17658 13375 17766 13485 4 gnd
port 517 nsew
rlabel metal2 s 15930 15525 16038 15601 4 gnd
port 517 nsew
rlabel metal2 s 18426 17325 18534 17435 4 gnd
port 517 nsew
rlabel metal2 s 186 9679 294 9755 4 gnd
port 517 nsew
rlabel metal2 s 186 18115 294 18225 4 gnd
port 517 nsew
rlabel metal2 s 2202 19949 2310 20025 4 gnd
port 517 nsew
rlabel metal2 s 18906 19159 19014 19235 4 gnd
port 517 nsew
rlabel metal2 s 3450 21275 3558 21385 4 gnd
port 517 nsew
rlabel metal2 s 15162 19695 15270 19805 4 gnd
port 517 nsew
rlabel metal2 s 5946 9995 6054 10071 4 gnd
port 517 nsew
rlabel metal2 s 11418 23645 11526 23755 4 gnd
port 517 nsew
rlabel metal2 s 12186 24689 12294 24765 4 gnd
port 517 nsew
rlabel metal2 s 1434 22635 1542 22711 4 gnd
port 517 nsew
rlabel metal2 s 3930 515 4038 591 4 gnd
port 517 nsew
rlabel metal2 s 5178 17325 5286 17435 4 gnd
port 517 nsew
rlabel metal2 s 16410 2885 16518 2961 4 gnd
port 517 nsew
rlabel metal2 s 12666 9425 12774 9535 4 gnd
port 517 nsew
rlabel metal2 s 14682 23899 14790 23975 4 gnd
port 517 nsew
rlabel metal2 s 15162 6519 15270 6595 4 gnd
port 517 nsew
rlabel metal2 s 8442 22635 8550 22711 4 gnd
port 517 nsew
rlabel metal2 s 17178 14165 17286 14275 4 gnd
port 517 nsew
rlabel metal2 s 10170 7309 10278 7385 4 gnd
port 517 nsew
rlabel metal2 s 5946 5729 6054 5805 4 gnd
port 517 nsew
rlabel metal2 s 10170 10785 10278 10861 4 gnd
port 517 nsew
rlabel metal2 s 9690 2569 9798 2645 4 gnd
port 517 nsew
rlabel metal2 s 15162 22635 15270 22711 4 gnd
port 517 nsew
rlabel metal2 s 18906 22065 19014 22175 4 gnd
port 517 nsew
rlabel metal2 s 3450 20739 3558 20815 4 gnd
port 517 nsew
rlabel metal2 s 7194 2885 7302 2961 4 gnd
port 517 nsew
rlabel metal2 s 10170 23899 10278 23975 4 gnd
port 517 nsew
rlabel metal2 s 5178 11259 5286 11335 4 gnd
port 517 nsew
rlabel metal2 s 10938 1779 11046 1855 4 gnd
port 517 nsew
rlabel metal2 s 15162 6835 15270 6911 4 gnd
port 517 nsew
rlabel metal2 s 954 9205 1062 9281 4 gnd
port 517 nsew
rlabel metal2 s 15930 25225 16038 25335 4 gnd
port 517 nsew
rlabel metal2 s 186 10785 294 10861 4 gnd
port 517 nsew
rlabel metal2 s 3930 1305 4038 1381 4 gnd
port 517 nsew
rlabel metal2 s 5946 515 6054 591 4 gnd
port 517 nsew
rlabel metal2 s 10938 9425 11046 9535 4 gnd
port 517 nsew
rlabel metal2 s 8922 11795 9030 11905 4 gnd
port 517 nsew
rlabel metal2 s 3930 5255 4038 5331 4 gnd
port 517 nsew
rlabel metal2 s 9690 12049 9798 12125 4 gnd
port 517 nsew
rlabel metal2 s 10938 8635 11046 8745 4 gnd
port 517 nsew
rlabel metal2 s 11418 2095 11526 2171 4 gnd
port 517 nsew
rlabel metal2 s 954 12839 1062 12915 4 gnd
port 517 nsew
rlabel metal2 s 7194 11795 7302 11905 4 gnd
port 517 nsew
rlabel metal2 s 9690 11795 9798 11905 4 gnd
port 517 nsew
rlabel metal2 s 18906 2885 19014 2961 4 gnd
port 517 nsew
rlabel metal2 s 16410 14735 16518 14811 4 gnd
port 517 nsew
rlabel metal2 s 8922 1525 9030 1635 4 gnd
port 517 nsew
rlabel metal2 s 186 21055 294 21131 4 gnd
port 517 nsew
rlabel metal2 s 12186 4465 12294 4541 4 gnd
port 517 nsew
rlabel metal2 s 1434 1779 1542 1855 4 gnd
port 517 nsew
rlabel metal2 s 3450 3359 3558 3435 4 gnd
port 517 nsew
rlabel metal2 s 954 21529 1062 21605 4 gnd
port 517 nsew
rlabel metal2 s 13914 15525 14022 15601 4 gnd
port 517 nsew
rlabel metal2 s 12666 4685 12774 4795 4 gnd
port 517 nsew
rlabel metal2 s 17178 19159 17286 19235 4 gnd
port 517 nsew
rlabel metal2 s 186 19475 294 19551 4 gnd
port 517 nsew
rlabel metal2 s 3450 12049 3558 12125 4 gnd
port 517 nsew
rlabel metal2 s 6426 1779 6534 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 1779 7782 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 4149 7782 4225 4 gnd
port 517 nsew
rlabel metal2 s 9690 13629 9798 13705 4 gnd
port 517 nsew
rlabel metal2 s 17658 6265 17766 6375 4 gnd
port 517 nsew
rlabel metal2 s 1434 8635 1542 8745 4 gnd
port 517 nsew
rlabel metal2 s 12666 15209 12774 15285 4 gnd
port 517 nsew
rlabel metal2 s 10170 6045 10278 6121 4 gnd
port 517 nsew
rlabel metal2 s 954 2095 1062 2171 4 gnd
port 517 nsew
rlabel metal2 s 18906 14955 19014 15065 4 gnd
port 517 nsew
rlabel metal2 s 11418 735 11526 845 4 gnd
port 517 nsew
rlabel metal2 s 1434 23425 1542 23501 4 gnd
port 517 nsew
rlabel metal2 s 15162 989 15270 1065 4 gnd
port 517 nsew
rlabel metal2 s 15162 17105 15270 17181 4 gnd
port 517 nsew
rlabel metal2 s 19674 12585 19782 12695 4 gnd
port 517 nsew
rlabel metal2 s 18426 6045 18534 6121 4 gnd
port 517 nsew
rlabel metal2 s 6426 17325 6534 17435 4 gnd
port 517 nsew
rlabel metal2 s 2682 14165 2790 14275 4 gnd
port 517 nsew
rlabel metal2 s 8442 3105 8550 3215 4 gnd
port 517 nsew
rlabel metal2 s 3930 22319 4038 22395 4 gnd
port 517 nsew
rlabel metal2 s 2682 8415 2790 8491 4 gnd
port 517 nsew
rlabel metal2 s 3930 25005 4038 25081 4 gnd
port 517 nsew
rlabel metal2 s 15930 515 16038 591 4 gnd
port 517 nsew
rlabel metal2 s 12186 6519 12294 6595 4 gnd
port 517 nsew
rlabel metal2 s 12186 15525 12294 15601 4 gnd
port 517 nsew
rlabel metal2 s 9690 14165 9798 14275 4 gnd
port 517 nsew
rlabel metal2 s 18906 9995 19014 10071 4 gnd
port 517 nsew
rlabel metal2 s 19674 735 19782 845 4 gnd
port 517 nsew
rlabel metal2 s 3930 1779 4038 1855 4 gnd
port 517 nsew
rlabel metal2 s 10938 12839 11046 12915 4 gnd
port 517 nsew
rlabel metal2 s 11418 10469 11526 10545 4 gnd
port 517 nsew
rlabel metal2 s 12666 11795 12774 11905 4 gnd
port 517 nsew
rlabel metal2 s 5178 21275 5286 21385 4 gnd
port 517 nsew
rlabel metal2 s 11418 21845 11526 21921 4 gnd
port 517 nsew
rlabel metal2 s 17658 21845 17766 21921 4 gnd
port 517 nsew
rlabel metal2 s 2682 17579 2790 17655 4 gnd
port 517 nsew
rlabel metal2 s 7194 9205 7302 9281 4 gnd
port 517 nsew
rlabel metal2 s 8922 12049 9030 12125 4 gnd
port 517 nsew
rlabel metal2 s 3450 1305 3558 1381 4 gnd
port 517 nsew
rlabel metal2 s 16410 735 16518 845 4 gnd
port 517 nsew
rlabel metal2 s 17178 23425 17286 23501 4 gnd
port 517 nsew
rlabel metal2 s 12666 15525 12774 15601 4 gnd
port 517 nsew
rlabel metal2 s 15930 23645 16038 23755 4 gnd
port 517 nsew
rlabel metal2 s 5946 16315 6054 16391 4 gnd
port 517 nsew
rlabel metal2 s 14682 18115 14790 18225 4 gnd
port 517 nsew
rlabel metal2 s 2682 19695 2790 19805 4 gnd
port 517 nsew
rlabel metal2 s 13434 5255 13542 5331 4 gnd
port 517 nsew
rlabel metal2 s 15930 1779 16038 1855 4 gnd
port 517 nsew
rlabel metal2 s 19674 19475 19782 19551 4 gnd
port 517 nsew
rlabel metal2 s 2202 11259 2310 11335 4 gnd
port 517 nsew
rlabel metal2 s 12666 19475 12774 19551 4 gnd
port 517 nsew
rlabel metal2 s 15162 19159 15270 19235 4 gnd
port 517 nsew
rlabel metal2 s 6426 12049 6534 12125 4 gnd
port 517 nsew
rlabel metal2 s 15930 17325 16038 17435 4 gnd
port 517 nsew
rlabel metal2 s 13434 15525 13542 15601 4 gnd
port 517 nsew
rlabel metal2 s 2202 5475 2310 5585 4 gnd
port 517 nsew
rlabel metal2 s 6426 7625 6534 7701 4 gnd
port 517 nsew
rlabel metal2 s 6426 1305 6534 1381 4 gnd
port 517 nsew
rlabel metal2 s 15930 4685 16038 4795 4 gnd
port 517 nsew
rlabel metal2 s 4698 13945 4806 14021 4 gnd
port 517 nsew
rlabel metal2 s 10170 9425 10278 9535 4 gnd
port 517 nsew
rlabel metal2 s 2202 1525 2310 1635 4 gnd
port 517 nsew
rlabel metal2 s 9690 8889 9798 8965 4 gnd
port 517 nsew
rlabel metal2 s 2682 19949 2790 20025 4 gnd
port 517 nsew
rlabel metal2 s 3930 14419 4038 14495 4 gnd
port 517 nsew
rlabel metal2 s 7194 21845 7302 21921 4 gnd
port 517 nsew
rlabel metal2 s 186 4149 294 4225 4 gnd
port 517 nsew
rlabel metal2 s 14682 15745 14790 15855 4 gnd
port 517 nsew
rlabel metal2 s 12666 -55 12774 55 4 gnd
port 517 nsew
rlabel metal2 s 14682 12049 14790 12125 4 gnd
port 517 nsew
rlabel metal2 s 17658 13155 17766 13231 4 gnd
port 517 nsew
rlabel metal2 s 4698 735 4806 845 4 gnd
port 517 nsew
rlabel metal2 s 8922 10215 9030 10325 4 gnd
port 517 nsew
rlabel metal2 s 18426 1305 18534 1381 4 gnd
port 517 nsew
rlabel metal2 s 13914 4939 14022 5015 4 gnd
port 517 nsew
rlabel metal2 s 3930 4149 4038 4225 4 gnd
port 517 nsew
rlabel metal2 s 9690 12365 9798 12441 4 gnd
port 517 nsew
rlabel metal2 s 12186 9205 12294 9281 4 gnd
port 517 nsew
rlabel metal2 s 186 20485 294 20595 4 gnd
port 517 nsew
rlabel metal2 s 5946 17579 6054 17655 4 gnd
port 517 nsew
rlabel metal2 s 12666 19159 12774 19235 4 gnd
port 517 nsew
rlabel metal2 s 12186 12049 12294 12125 4 gnd
port 517 nsew
rlabel metal2 s 10170 21055 10278 21131 4 gnd
port 517 nsew
rlabel metal2 s 5178 24435 5286 24545 4 gnd
port 517 nsew
rlabel metal2 s 11418 989 11526 1065 4 gnd
port 517 nsew
rlabel metal2 s 3450 3675 3558 3751 4 gnd
port 517 nsew
rlabel metal2 s 16410 8415 16518 8491 4 gnd
port 517 nsew
rlabel metal2 s 5178 4149 5286 4225 4 gnd
port 517 nsew
rlabel metal2 s 1434 14955 1542 15065 4 gnd
port 517 nsew
rlabel metal2 s 1434 17105 1542 17181 4 gnd
port 517 nsew
rlabel metal2 s 5178 23425 5286 23501 4 gnd
port 517 nsew
rlabel metal2 s 954 11575 1062 11651 4 gnd
port 517 nsew
rlabel metal2 s 954 8889 1062 8965 4 gnd
port 517 nsew
rlabel metal2 s 1434 9205 1542 9281 4 gnd
port 517 nsew
rlabel metal2 s 3450 4685 3558 4795 4 gnd
port 517 nsew
rlabel metal2 s 7674 12585 7782 12695 4 gnd
port 517 nsew
rlabel metal2 s 8442 11259 8550 11335 4 gnd
port 517 nsew
rlabel metal2 s 5946 10785 6054 10861 4 gnd
port 517 nsew
rlabel metal2 s 8442 8635 8550 8745 4 gnd
port 517 nsew
rlabel metal2 s 954 22319 1062 22395 4 gnd
port 517 nsew
rlabel metal2 s 8922 23425 9030 23501 4 gnd
port 517 nsew
rlabel metal2 s 11418 8635 11526 8745 4 gnd
port 517 nsew
rlabel metal2 s 13434 10469 13542 10545 4 gnd
port 517 nsew
rlabel metal2 s 186 13375 294 13485 4 gnd
port 517 nsew
rlabel metal2 s 10938 13155 11046 13231 4 gnd
port 517 nsew
rlabel metal2 s 11418 9205 11526 9281 4 gnd
port 517 nsew
rlabel metal2 s 17658 18115 17766 18225 4 gnd
port 517 nsew
rlabel metal2 s 7194 8889 7302 8965 4 gnd
port 517 nsew
rlabel metal2 s 12666 16535 12774 16645 4 gnd
port 517 nsew
rlabel metal2 s 2682 16535 2790 16645 4 gnd
port 517 nsew
rlabel metal2 s 5946 13629 6054 13705 4 gnd
port 517 nsew
rlabel metal2 s 12186 15999 12294 16075 4 gnd
port 517 nsew
rlabel metal2 s 5178 6265 5286 6375 4 gnd
port 517 nsew
rlabel metal2 s 14682 5729 14790 5805 4 gnd
port 517 nsew
rlabel metal2 s 7194 9425 7302 9535 4 gnd
port 517 nsew
rlabel metal2 s 19674 1305 19782 1381 4 gnd
port 517 nsew
rlabel metal2 s 12666 13375 12774 13485 4 gnd
port 517 nsew
rlabel metal2 s 18426 21529 18534 21605 4 gnd
port 517 nsew
rlabel metal2 s 12186 4149 12294 4225 4 gnd
port 517 nsew
rlabel metal2 s 12186 15745 12294 15855 4 gnd
port 517 nsew
rlabel metal2 s 3930 4465 4038 4541 4 gnd
port 517 nsew
rlabel metal2 s 15930 23899 16038 23975 4 gnd
port 517 nsew
rlabel metal2 s 9690 7055 9798 7165 4 gnd
port 517 nsew
rlabel metal2 s 9690 20739 9798 20815 4 gnd
port 517 nsew
rlabel metal2 s 15162 16535 15270 16645 4 gnd
port 517 nsew
rlabel metal2 s 17178 18115 17286 18225 4 gnd
port 517 nsew
rlabel metal2 s 12666 1305 12774 1381 4 gnd
port 517 nsew
rlabel metal2 s 10170 1779 10278 1855 4 gnd
port 517 nsew
rlabel metal2 s 3930 14165 4038 14275 4 gnd
port 517 nsew
rlabel metal2 s 19674 19695 19782 19805 4 gnd
port 517 nsew
rlabel metal2 s 18906 16535 19014 16645 4 gnd
port 517 nsew
rlabel metal2 s 3450 4939 3558 5015 4 gnd
port 517 nsew
rlabel metal2 s 954 7625 1062 7701 4 gnd
port 517 nsew
rlabel metal2 s 13914 8889 14022 8965 4 gnd
port 517 nsew
rlabel metal2 s 2682 17895 2790 17971 4 gnd
port 517 nsew
rlabel metal2 s 6426 11795 6534 11905 4 gnd
port 517 nsew
rlabel metal2 s 8922 17579 9030 17655 4 gnd
port 517 nsew
rlabel metal2 s 12666 1779 12774 1855 4 gnd
port 517 nsew
rlabel metal2 s 8922 7625 9030 7701 4 gnd
port 517 nsew
rlabel metal2 s 13434 2095 13542 2171 4 gnd
port 517 nsew
rlabel metal2 s 1434 19695 1542 19805 4 gnd
port 517 nsew
rlabel metal2 s 2682 15999 2790 16075 4 gnd
port 517 nsew
rlabel metal2 s 14682 20485 14790 20595 4 gnd
port 517 nsew
rlabel metal2 s 19674 7309 19782 7385 4 gnd
port 517 nsew
rlabel metal2 s 186 10215 294 10325 4 gnd
port 517 nsew
rlabel metal2 s 19674 16535 19782 16645 4 gnd
port 517 nsew
rlabel metal2 s 3930 7845 4038 7955 4 gnd
port 517 nsew
rlabel metal2 s 10938 4149 11046 4225 4 gnd
port 517 nsew
rlabel metal2 s 14682 10215 14790 10325 4 gnd
port 517 nsew
rlabel metal2 s 186 11795 294 11905 4 gnd
port 517 nsew
rlabel metal2 s 2202 2885 2310 2961 4 gnd
port 517 nsew
rlabel metal2 s 5178 18685 5286 18761 4 gnd
port 517 nsew
rlabel metal2 s 13434 24215 13542 24291 4 gnd
port 517 nsew
rlabel metal2 s 15930 6265 16038 6375 4 gnd
port 517 nsew
rlabel metal2 s 16410 12049 16518 12125 4 gnd
port 517 nsew
rlabel metal2 s 8442 8415 8550 8491 4 gnd
port 517 nsew
rlabel metal2 s 16410 21055 16518 21131 4 gnd
port 517 nsew
rlabel metal2 s 3450 199 3558 275 4 gnd
port 517 nsew
rlabel metal2 s 12186 4939 12294 5015 4 gnd
port 517 nsew
rlabel metal2 s 3450 16315 3558 16391 4 gnd
port 517 nsew
rlabel metal2 s 11418 18905 11526 19015 4 gnd
port 517 nsew
rlabel metal2 s 12186 13375 12294 13485 4 gnd
port 517 nsew
rlabel metal2 s 13914 17895 14022 17971 4 gnd
port 517 nsew
rlabel metal2 s 18906 4465 19014 4541 4 gnd
port 517 nsew
rlabel metal2 s 18906 20265 19014 20341 4 gnd
port 517 nsew
rlabel metal2 s 3930 17105 4038 17181 4 gnd
port 517 nsew
rlabel metal2 s 15162 14735 15270 14811 4 gnd
port 517 nsew
rlabel metal2 s 11418 6835 11526 6911 4 gnd
port 517 nsew
rlabel metal2 s 10938 735 11046 845 4 gnd
port 517 nsew
rlabel metal2 s 11418 14419 11526 14495 4 gnd
port 517 nsew
rlabel metal2 s 13914 23899 14022 23975 4 gnd
port 517 nsew
rlabel metal2 s 19674 15745 19782 15855 4 gnd
port 517 nsew
rlabel metal2 s 1434 2095 1542 2171 4 gnd
port 517 nsew
rlabel metal2 s 12186 9995 12294 10071 4 gnd
port 517 nsew
rlabel metal2 s 7674 4465 7782 4541 4 gnd
port 517 nsew
rlabel metal2 s 10938 15745 11046 15855 4 gnd
port 517 nsew
rlabel metal2 s 11418 16315 11526 16391 4 gnd
port 517 nsew
rlabel metal2 s 6426 14955 6534 15065 4 gnd
port 517 nsew
rlabel metal2 s 10170 15745 10278 15855 4 gnd
port 517 nsew
rlabel metal2 s 14682 18905 14790 19015 4 gnd
port 517 nsew
rlabel metal2 s 8922 22855 9030 22965 4 gnd
port 517 nsew
rlabel metal2 s 17658 9679 17766 9755 4 gnd
port 517 nsew
rlabel metal2 s 17658 20485 17766 20595 4 gnd
port 517 nsew
rlabel metal2 s 17658 12365 17766 12441 4 gnd
port 517 nsew
rlabel metal2 s 5178 2885 5286 2961 4 gnd
port 517 nsew
rlabel metal2 s 17658 11795 17766 11905 4 gnd
port 517 nsew
rlabel metal2 s 2202 9425 2310 9535 4 gnd
port 517 nsew
rlabel metal2 s 954 11005 1062 11115 4 gnd
port 517 nsew
rlabel metal2 s 17178 3105 17286 3215 4 gnd
port 517 nsew
rlabel metal2 s 3930 9425 4038 9535 4 gnd
port 517 nsew
rlabel metal2 s 7674 14955 7782 15065 4 gnd
port 517 nsew
rlabel metal2 s 7674 3675 7782 3751 4 gnd
port 517 nsew
rlabel metal2 s 8442 17105 8550 17181 4 gnd
port 517 nsew
rlabel metal2 s 17658 24689 17766 24765 4 gnd
port 517 nsew
rlabel metal2 s 12186 989 12294 1065 4 gnd
port 517 nsew
rlabel metal2 s 18426 4149 18534 4225 4 gnd
port 517 nsew
rlabel metal2 s 6426 20739 6534 20815 4 gnd
port 517 nsew
rlabel metal2 s 16410 1305 16518 1381 4 gnd
port 517 nsew
rlabel metal2 s 16410 21529 16518 21605 4 gnd
port 517 nsew
rlabel metal2 s 8922 3675 9030 3751 4 gnd
port 517 nsew
rlabel metal2 s 12666 22319 12774 22395 4 gnd
port 517 nsew
rlabel metal2 s 18906 12365 19014 12441 4 gnd
port 517 nsew
rlabel metal2 s 7194 20265 7302 20341 4 gnd
port 517 nsew
rlabel metal2 s 8922 21845 9030 21921 4 gnd
port 517 nsew
rlabel metal2 s 8442 23645 8550 23755 4 gnd
port 517 nsew
rlabel metal2 s 9690 23109 9798 23185 4 gnd
port 517 nsew
rlabel metal2 s 17658 23899 17766 23975 4 gnd
port 517 nsew
rlabel metal2 s 186 12365 294 12441 4 gnd
port 517 nsew
rlabel metal2 s 10938 6835 11046 6911 4 gnd
port 517 nsew
rlabel metal2 s 16410 15525 16518 15601 4 gnd
port 517 nsew
rlabel metal2 s 5946 18905 6054 19015 4 gnd
port 517 nsew
rlabel metal2 s 18426 7309 18534 7385 4 gnd
port 517 nsew
rlabel metal2 s 4698 3105 4806 3215 4 gnd
port 517 nsew
rlabel metal2 s 15162 18115 15270 18225 4 gnd
port 517 nsew
rlabel metal2 s 3450 6519 3558 6595 4 gnd
port 517 nsew
rlabel metal2 s 13914 24435 14022 24545 4 gnd
port 517 nsew
rlabel metal2 s 10170 989 10278 1065 4 gnd
port 517 nsew
rlabel metal2 s 8922 4685 9030 4795 4 gnd
port 517 nsew
rlabel metal2 s 18906 2569 19014 2645 4 gnd
port 517 nsew
rlabel metal2 s 18906 17579 19014 17655 4 gnd
port 517 nsew
rlabel metal2 s 11418 3359 11526 3435 4 gnd
port 517 nsew
rlabel metal2 s 6426 11005 6534 11115 4 gnd
port 517 nsew
rlabel metal2 s 5178 2095 5286 2171 4 gnd
port 517 nsew
rlabel metal2 s 3930 25225 4038 25335 4 gnd
port 517 nsew
rlabel metal2 s 5946 13155 6054 13231 4 gnd
port 517 nsew
rlabel metal2 s 5946 3675 6054 3751 4 gnd
port 517 nsew
rlabel metal2 s 186 14955 294 15065 4 gnd
port 517 nsew
rlabel metal2 s 17178 12049 17286 12125 4 gnd
port 517 nsew
rlabel metal2 s 12666 25005 12774 25081 4 gnd
port 517 nsew
rlabel metal2 s 4698 19949 4806 20025 4 gnd
port 517 nsew
rlabel metal2 s 7674 22065 7782 22175 4 gnd
port 517 nsew
rlabel metal2 s 15930 9205 16038 9281 4 gnd
port 517 nsew
rlabel metal2 s 5946 3359 6054 3435 4 gnd
port 517 nsew
rlabel metal2 s 12666 3105 12774 3215 4 gnd
port 517 nsew
rlabel metal2 s 17658 17105 17766 17181 4 gnd
port 517 nsew
rlabel metal2 s 2202 20485 2310 20595 4 gnd
port 517 nsew
rlabel metal2 s 14682 19949 14790 20025 4 gnd
port 517 nsew
rlabel metal2 s 9690 4939 9798 5015 4 gnd
port 517 nsew
rlabel metal2 s 5178 11005 5286 11115 4 gnd
port 517 nsew
rlabel metal2 s 8442 11005 8550 11115 4 gnd
port 517 nsew
rlabel metal2 s 17178 4939 17286 5015 4 gnd
port 517 nsew
rlabel metal2 s 7194 16535 7302 16645 4 gnd
port 517 nsew
rlabel metal2 s 15930 2569 16038 2645 4 gnd
port 517 nsew
rlabel metal2 s 2682 -55 2790 55 4 gnd
port 517 nsew
rlabel metal2 s 15162 4149 15270 4225 4 gnd
port 517 nsew
rlabel metal2 s 10170 13375 10278 13485 4 gnd
port 517 nsew
rlabel metal2 s 1434 9995 1542 10071 4 gnd
port 517 nsew
rlabel metal2 s 2202 22635 2310 22711 4 gnd
port 517 nsew
rlabel metal2 s 12186 20739 12294 20815 4 gnd
port 517 nsew
rlabel metal2 s 14682 15209 14790 15285 4 gnd
port 517 nsew
rlabel metal2 s 11418 24689 11526 24765 4 gnd
port 517 nsew
rlabel metal2 s 16410 14955 16518 15065 4 gnd
port 517 nsew
rlabel metal2 s 10170 12839 10278 12915 4 gnd
port 517 nsew
rlabel metal2 s 15930 24215 16038 24291 4 gnd
port 517 nsew
rlabel metal2 s 3450 18369 3558 18445 4 gnd
port 517 nsew
rlabel metal2 s 2202 18369 2310 18445 4 gnd
port 517 nsew
rlabel metal2 s 12666 23645 12774 23755 4 gnd
port 517 nsew
rlabel metal2 s 10938 23109 11046 23185 4 gnd
port 517 nsew
rlabel metal2 s 6426 15999 6534 16075 4 gnd
port 517 nsew
rlabel metal2 s 3450 25225 3558 25335 4 gnd
port 517 nsew
rlabel metal2 s 186 9995 294 10071 4 gnd
port 517 nsew
rlabel metal2 s 1434 24215 1542 24291 4 gnd
port 517 nsew
rlabel metal2 s 3450 18115 3558 18225 4 gnd
port 517 nsew
rlabel metal2 s 18426 24689 18534 24765 4 gnd
port 517 nsew
rlabel metal2 s 12186 -55 12294 55 4 gnd
port 517 nsew
rlabel metal2 s 10170 4149 10278 4225 4 gnd
port 517 nsew
rlabel metal2 s 954 5475 1062 5585 4 gnd
port 517 nsew
rlabel metal2 s 2682 24689 2790 24765 4 gnd
port 517 nsew
rlabel metal2 s 16410 3895 16518 4005 4 gnd
port 517 nsew
rlabel metal2 s 17178 6045 17286 6121 4 gnd
port 517 nsew
rlabel metal2 s 7674 2315 7782 2425 4 gnd
port 517 nsew
rlabel metal2 s 17658 2095 17766 2171 4 gnd
port 517 nsew
rlabel metal2 s 3930 15999 4038 16075 4 gnd
port 517 nsew
rlabel metal2 s 5946 15999 6054 16075 4 gnd
port 517 nsew
rlabel metal2 s 8922 8889 9030 8965 4 gnd
port 517 nsew
rlabel metal2 s 4698 4685 4806 4795 4 gnd
port 517 nsew
rlabel metal2 s 5946 4685 6054 4795 4 gnd
port 517 nsew
rlabel metal2 s 18426 8889 18534 8965 4 gnd
port 517 nsew
rlabel metal2 s 15930 4465 16038 4541 4 gnd
port 517 nsew
rlabel metal2 s 8922 17895 9030 17971 4 gnd
port 517 nsew
rlabel metal2 s 6426 7309 6534 7385 4 gnd
port 517 nsew
rlabel metal2 s 8442 9679 8550 9755 4 gnd
port 517 nsew
rlabel metal2 s 3930 13375 4038 13485 4 gnd
port 517 nsew
rlabel metal2 s 954 10215 1062 10325 4 gnd
port 517 nsew
rlabel metal2 s 10170 23109 10278 23185 4 gnd
port 517 nsew
rlabel metal2 s 10170 15525 10278 15601 4 gnd
port 517 nsew
rlabel metal2 s 11418 5475 11526 5585 4 gnd
port 517 nsew
rlabel metal2 s 6426 2885 6534 2961 4 gnd
port 517 nsew
rlabel metal2 s 5178 6045 5286 6121 4 gnd
port 517 nsew
rlabel metal2 s 3450 19695 3558 19805 4 gnd
port 517 nsew
rlabel metal2 s 10170 24215 10278 24291 4 gnd
port 517 nsew
rlabel metal2 s 3930 10469 4038 10545 4 gnd
port 517 nsew
rlabel metal2 s 18906 14419 19014 14495 4 gnd
port 517 nsew
rlabel metal2 s 14682 3359 14790 3435 4 gnd
port 517 nsew
rlabel metal2 s 17658 5729 17766 5805 4 gnd
port 517 nsew
rlabel metal2 s 18906 199 19014 275 4 gnd
port 517 nsew
rlabel metal2 s 954 17105 1062 17181 4 gnd
port 517 nsew
rlabel metal2 s 9690 3359 9798 3435 4 gnd
port 517 nsew
rlabel metal2 s 10170 25005 10278 25081 4 gnd
port 517 nsew
rlabel metal2 s 17178 1525 17286 1635 4 gnd
port 517 nsew
rlabel metal2 s 19674 18369 19782 18445 4 gnd
port 517 nsew
rlabel metal2 s 17658 10469 17766 10545 4 gnd
port 517 nsew
rlabel metal2 s 12666 7055 12774 7165 4 gnd
port 517 nsew
rlabel metal2 s 18906 18369 19014 18445 4 gnd
port 517 nsew
rlabel metal2 s 9690 23899 9798 23975 4 gnd
port 517 nsew
rlabel metal2 s 954 1525 1062 1635 4 gnd
port 517 nsew
rlabel metal2 s 12666 515 12774 591 4 gnd
port 517 nsew
rlabel metal2 s 13914 2315 14022 2425 4 gnd
port 517 nsew
rlabel metal2 s 11418 2885 11526 2961 4 gnd
port 517 nsew
rlabel metal2 s 186 11005 294 11115 4 gnd
port 517 nsew
rlabel metal2 s 2202 2095 2310 2171 4 gnd
port 517 nsew
rlabel metal2 s 15930 18369 16038 18445 4 gnd
port 517 nsew
rlabel metal2 s 2682 25225 2790 25335 4 gnd
port 517 nsew
rlabel metal2 s 15162 20265 15270 20341 4 gnd
port 517 nsew
rlabel metal2 s 14682 16315 14790 16391 4 gnd
port 517 nsew
rlabel metal2 s 186 10469 294 10545 4 gnd
port 517 nsew
rlabel metal2 s 3450 1525 3558 1635 4 gnd
port 517 nsew
rlabel metal2 s 19674 21055 19782 21131 4 gnd
port 517 nsew
rlabel metal2 s 13914 5255 14022 5331 4 gnd
port 517 nsew
rlabel metal2 s 14682 10785 14790 10861 4 gnd
port 517 nsew
rlabel metal2 s 12666 11005 12774 11115 4 gnd
port 517 nsew
rlabel metal2 s 18426 7055 18534 7165 4 gnd
port 517 nsew
rlabel metal2 s 7194 4685 7302 4795 4 gnd
port 517 nsew
rlabel metal2 s 7674 22855 7782 22965 4 gnd
port 517 nsew
rlabel metal2 s 3450 22319 3558 22395 4 gnd
port 517 nsew
rlabel metal2 s 2682 2885 2790 2961 4 gnd
port 517 nsew
rlabel metal2 s 12186 3359 12294 3435 4 gnd
port 517 nsew
rlabel metal2 s 18426 5255 18534 5331 4 gnd
port 517 nsew
rlabel metal2 s 16410 9205 16518 9281 4 gnd
port 517 nsew
rlabel metal2 s 17178 -55 17286 55 4 gnd
port 517 nsew
rlabel metal2 s 13914 11575 14022 11651 4 gnd
port 517 nsew
rlabel metal2 s 18906 21055 19014 21131 4 gnd
port 517 nsew
rlabel metal2 s 5178 11795 5286 11905 4 gnd
port 517 nsew
rlabel metal2 s 8442 5475 8550 5585 4 gnd
port 517 nsew
rlabel metal2 s 5946 6265 6054 6375 4 gnd
port 517 nsew
rlabel metal2 s 11418 3675 11526 3751 4 gnd
port 517 nsew
rlabel metal2 s 16410 14419 16518 14495 4 gnd
port 517 nsew
rlabel metal2 s 18426 7845 18534 7955 4 gnd
port 517 nsew
rlabel metal2 s 954 11259 1062 11335 4 gnd
port 517 nsew
rlabel metal2 s 19674 3105 19782 3215 4 gnd
port 517 nsew
rlabel metal2 s 1434 9679 1542 9755 4 gnd
port 517 nsew
rlabel metal2 s 15162 2095 15270 2171 4 gnd
port 517 nsew
rlabel metal2 s 5946 15525 6054 15601 4 gnd
port 517 nsew
rlabel metal2 s 14682 4465 14790 4541 4 gnd
port 517 nsew
rlabel metal2 s 10170 15999 10278 16075 4 gnd
port 517 nsew
rlabel metal2 s 9690 24215 9798 24291 4 gnd
port 517 nsew
rlabel metal2 s 6426 4465 6534 4541 4 gnd
port 517 nsew
rlabel metal2 s 10938 11795 11046 11905 4 gnd
port 517 nsew
rlabel metal2 s 2682 8635 2790 8745 4 gnd
port 517 nsew
rlabel metal2 s 18426 1779 18534 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 20485 7782 20595 4 gnd
port 517 nsew
rlabel metal2 s 10938 21845 11046 21921 4 gnd
port 517 nsew
rlabel metal2 s 1434 9425 1542 9535 4 gnd
port 517 nsew
rlabel metal2 s 10938 17579 11046 17655 4 gnd
port 517 nsew
rlabel metal2 s 186 24215 294 24291 4 gnd
port 517 nsew
rlabel metal2 s 5946 19159 6054 19235 4 gnd
port 517 nsew
rlabel metal2 s 17658 8635 17766 8745 4 gnd
port 517 nsew
rlabel metal2 s 11418 4465 11526 4541 4 gnd
port 517 nsew
rlabel metal2 s 954 12049 1062 12125 4 gnd
port 517 nsew
rlabel metal2 s 18906 7055 19014 7165 4 gnd
port 517 nsew
rlabel metal2 s 2202 7845 2310 7955 4 gnd
port 517 nsew
rlabel metal2 s 3930 21275 4038 21385 4 gnd
port 517 nsew
rlabel metal2 s 15162 24435 15270 24545 4 gnd
port 517 nsew
rlabel metal2 s 16410 7625 16518 7701 4 gnd
port 517 nsew
rlabel metal2 s 12186 18115 12294 18225 4 gnd
port 517 nsew
rlabel metal2 s 18906 13629 19014 13705 4 gnd
port 517 nsew
rlabel metal2 s 19674 515 19782 591 4 gnd
port 517 nsew
rlabel metal2 s 5178 23109 5286 23185 4 gnd
port 517 nsew
rlabel metal2 s 12186 1779 12294 1855 4 gnd
port 517 nsew
rlabel metal2 s 3930 13155 4038 13231 4 gnd
port 517 nsew
rlabel metal2 s 10170 7625 10278 7701 4 gnd
port 517 nsew
rlabel metal2 s 9690 22855 9798 22965 4 gnd
port 517 nsew
rlabel metal2 s 4698 8099 4806 8175 4 gnd
port 517 nsew
rlabel metal2 s 8442 4685 8550 4795 4 gnd
port 517 nsew
rlabel metal2 s 1434 19949 1542 20025 4 gnd
port 517 nsew
rlabel metal2 s 18426 199 18534 275 4 gnd
port 517 nsew
rlabel metal2 s 11418 4149 11526 4225 4 gnd
port 517 nsew
rlabel metal2 s 2202 1305 2310 1381 4 gnd
port 517 nsew
rlabel metal2 s 9690 11005 9798 11115 4 gnd
port 517 nsew
rlabel metal2 s 11418 22635 11526 22711 4 gnd
port 517 nsew
rlabel metal2 s 16410 1779 16518 1855 4 gnd
port 517 nsew
rlabel metal2 s 12666 2315 12774 2425 4 gnd
port 517 nsew
rlabel metal2 s 3450 15525 3558 15601 4 gnd
port 517 nsew
rlabel metal2 s 17178 22065 17286 22175 4 gnd
port 517 nsew
rlabel metal2 s 8922 1779 9030 1855 4 gnd
port 517 nsew
rlabel metal2 s 186 17579 294 17655 4 gnd
port 517 nsew
rlabel metal2 s 14682 22065 14790 22175 4 gnd
port 517 nsew
rlabel metal2 s 2202 13629 2310 13705 4 gnd
port 517 nsew
rlabel metal2 s 7194 11259 7302 11335 4 gnd
port 517 nsew
rlabel metal2 s 8922 22319 9030 22395 4 gnd
port 517 nsew
rlabel metal2 s 8442 22855 8550 22965 4 gnd
port 517 nsew
rlabel metal2 s 18906 8415 19014 8491 4 gnd
port 517 nsew
rlabel metal2 s 15930 10215 16038 10325 4 gnd
port 517 nsew
rlabel metal2 s 10170 3675 10278 3751 4 gnd
port 517 nsew
rlabel metal2 s 13914 7055 14022 7165 4 gnd
port 517 nsew
rlabel metal2 s 18906 11795 19014 11905 4 gnd
port 517 nsew
rlabel metal2 s 19674 22065 19782 22175 4 gnd
port 517 nsew
rlabel metal2 s 2202 22065 2310 22175 4 gnd
port 517 nsew
rlabel metal2 s 13434 22319 13542 22395 4 gnd
port 517 nsew
rlabel metal2 s 7194 3105 7302 3215 4 gnd
port 517 nsew
rlabel metal2 s 3450 515 3558 591 4 gnd
port 517 nsew
rlabel metal2 s 15930 17895 16038 17971 4 gnd
port 517 nsew
rlabel metal2 s 8442 5729 8550 5805 4 gnd
port 517 nsew
rlabel metal2 s 7194 989 7302 1065 4 gnd
port 517 nsew
rlabel metal2 s 12186 11795 12294 11905 4 gnd
port 517 nsew
rlabel metal2 s 11418 23425 11526 23501 4 gnd
port 517 nsew
rlabel metal2 s 16410 17325 16518 17435 4 gnd
port 517 nsew
rlabel metal2 s 18426 18905 18534 19015 4 gnd
port 517 nsew
rlabel metal2 s 8442 11575 8550 11651 4 gnd
port 517 nsew
rlabel metal2 s 19674 17105 19782 17181 4 gnd
port 517 nsew
rlabel metal2 s 8922 5729 9030 5805 4 gnd
port 517 nsew
rlabel metal2 s 5178 10469 5286 10545 4 gnd
port 517 nsew
rlabel metal2 s 954 15209 1062 15285 4 gnd
port 517 nsew
rlabel metal2 s 16410 13375 16518 13485 4 gnd
port 517 nsew
rlabel metal2 s 9690 20485 9798 20595 4 gnd
port 517 nsew
rlabel metal2 s 5946 17895 6054 17971 4 gnd
port 517 nsew
rlabel metal2 s 8922 10785 9030 10861 4 gnd
port 517 nsew
rlabel metal2 s 10938 3359 11046 3435 4 gnd
port 517 nsew
rlabel metal2 s 13434 15999 13542 16075 4 gnd
port 517 nsew
rlabel metal2 s 15162 10215 15270 10325 4 gnd
port 517 nsew
rlabel metal2 s 14682 2885 14790 2961 4 gnd
port 517 nsew
rlabel metal2 s 18906 2315 19014 2425 4 gnd
port 517 nsew
rlabel metal2 s 12186 21275 12294 21385 4 gnd
port 517 nsew
rlabel metal2 s 4698 13375 4806 13485 4 gnd
port 517 nsew
rlabel metal2 s 3930 20739 4038 20815 4 gnd
port 517 nsew
rlabel metal2 s 2202 2569 2310 2645 4 gnd
port 517 nsew
rlabel metal2 s 5946 25005 6054 25081 4 gnd
port 517 nsew
rlabel metal2 s 7674 9679 7782 9755 4 gnd
port 517 nsew
rlabel metal2 s 6426 18905 6534 19015 4 gnd
port 517 nsew
rlabel metal2 s 8442 6045 8550 6121 4 gnd
port 517 nsew
rlabel metal2 s 10938 16789 11046 16865 4 gnd
port 517 nsew
rlabel metal2 s 17178 15209 17286 15285 4 gnd
port 517 nsew
rlabel metal2 s 15930 9425 16038 9535 4 gnd
port 517 nsew
rlabel metal2 s 11418 3895 11526 4005 4 gnd
port 517 nsew
rlabel metal2 s 3930 19695 4038 19805 4 gnd
port 517 nsew
rlabel metal2 s 5178 3359 5286 3435 4 gnd
port 517 nsew
rlabel metal2 s 954 1779 1062 1855 4 gnd
port 517 nsew
rlabel metal2 s 6426 7055 6534 7165 4 gnd
port 517 nsew
rlabel metal2 s 18906 21845 19014 21921 4 gnd
port 517 nsew
rlabel metal2 s 7674 6519 7782 6595 4 gnd
port 517 nsew
rlabel metal2 s 16410 199 16518 275 4 gnd
port 517 nsew
rlabel metal2 s 12666 23899 12774 23975 4 gnd
port 517 nsew
rlabel metal2 s 6426 12365 6534 12441 4 gnd
port 517 nsew
rlabel metal2 s 8922 2095 9030 2171 4 gnd
port 517 nsew
rlabel metal2 s 11418 17325 11526 17435 4 gnd
port 517 nsew
rlabel metal2 s 16410 13945 16518 14021 4 gnd
port 517 nsew
rlabel metal2 s 1434 16789 1542 16865 4 gnd
port 517 nsew
rlabel metal2 s 954 20739 1062 20815 4 gnd
port 517 nsew
rlabel metal2 s 8442 515 8550 591 4 gnd
port 517 nsew
rlabel metal2 s 954 735 1062 845 4 gnd
port 517 nsew
rlabel metal2 s 12186 21055 12294 21131 4 gnd
port 517 nsew
rlabel metal2 s 17658 23425 17766 23501 4 gnd
port 517 nsew
rlabel metal2 s 10170 16315 10278 16391 4 gnd
port 517 nsew
rlabel metal2 s 8922 14955 9030 15065 4 gnd
port 517 nsew
rlabel metal2 s 7194 -55 7302 55 4 gnd
port 517 nsew
rlabel metal2 s 5946 1779 6054 1855 4 gnd
port 517 nsew
rlabel metal2 s 9690 8635 9798 8745 4 gnd
port 517 nsew
rlabel metal2 s 13434 8099 13542 8175 4 gnd
port 517 nsew
rlabel metal2 s 1434 7309 1542 7385 4 gnd
port 517 nsew
rlabel metal2 s 19674 7845 19782 7955 4 gnd
port 517 nsew
rlabel metal2 s 4698 15745 4806 15855 4 gnd
port 517 nsew
rlabel metal2 s 10938 17895 11046 17971 4 gnd
port 517 nsew
rlabel metal2 s 5178 7309 5286 7385 4 gnd
port 517 nsew
rlabel metal2 s 10938 10215 11046 10325 4 gnd
port 517 nsew
rlabel metal2 s 3930 19159 4038 19235 4 gnd
port 517 nsew
rlabel metal2 s 5178 17895 5286 17971 4 gnd
port 517 nsew
rlabel metal2 s 19674 6265 19782 6375 4 gnd
port 517 nsew
rlabel metal2 s 19674 25225 19782 25335 4 gnd
port 517 nsew
rlabel metal2 s 954 8415 1062 8491 4 gnd
port 517 nsew
rlabel metal2 s 10938 18905 11046 19015 4 gnd
port 517 nsew
rlabel metal2 s 2202 1779 2310 1855 4 gnd
port 517 nsew
rlabel metal2 s 10938 15525 11046 15601 4 gnd
port 517 nsew
rlabel metal2 s 13434 2885 13542 2961 4 gnd
port 517 nsew
rlabel metal2 s 19674 2095 19782 2171 4 gnd
port 517 nsew
rlabel metal2 s 1434 21275 1542 21385 4 gnd
port 517 nsew
rlabel metal2 s 17178 3675 17286 3751 4 gnd
port 517 nsew
rlabel metal2 s 8442 2315 8550 2425 4 gnd
port 517 nsew
rlabel metal2 s 17658 19475 17766 19551 4 gnd
port 517 nsew
rlabel metal2 s 17658 20739 17766 20815 4 gnd
port 517 nsew
rlabel metal2 s 10170 9995 10278 10071 4 gnd
port 517 nsew
rlabel metal2 s 6426 25225 6534 25335 4 gnd
port 517 nsew
rlabel metal2 s 2682 9205 2790 9281 4 gnd
port 517 nsew
rlabel metal2 s 6426 -55 6534 55 4 gnd
port 517 nsew
rlabel metal2 s 3450 13155 3558 13231 4 gnd
port 517 nsew
rlabel metal2 s 5178 25005 5286 25081 4 gnd
port 517 nsew
rlabel metal2 s 3930 23425 4038 23501 4 gnd
port 517 nsew
rlabel metal2 s 11418 14735 11526 14811 4 gnd
port 517 nsew
rlabel metal2 s 2202 8635 2310 8745 4 gnd
port 517 nsew
rlabel metal2 s 11418 17579 11526 17655 4 gnd
port 517 nsew
rlabel metal2 s 15930 20485 16038 20595 4 gnd
port 517 nsew
rlabel metal2 s 15930 2885 16038 2961 4 gnd
port 517 nsew
rlabel metal2 s 16410 5255 16518 5331 4 gnd
port 517 nsew
rlabel metal2 s 7674 15745 7782 15855 4 gnd
port 517 nsew
rlabel metal2 s 17178 20265 17286 20341 4 gnd
port 517 nsew
rlabel metal2 s 4698 8889 4806 8965 4 gnd
port 517 nsew
rlabel metal2 s 17178 7055 17286 7165 4 gnd
port 517 nsew
rlabel metal2 s 7674 5475 7782 5585 4 gnd
port 517 nsew
rlabel metal2 s 17658 735 17766 845 4 gnd
port 517 nsew
rlabel metal2 s 10170 10469 10278 10545 4 gnd
port 517 nsew
rlabel metal2 s 15930 -55 16038 55 4 gnd
port 517 nsew
rlabel metal2 s 954 9679 1062 9755 4 gnd
port 517 nsew
rlabel metal2 s 10170 20485 10278 20595 4 gnd
port 517 nsew
rlabel metal2 s 12186 16535 12294 16645 4 gnd
port 517 nsew
rlabel metal2 s 12666 22065 12774 22175 4 gnd
port 517 nsew
rlabel metal2 s 17178 15525 17286 15601 4 gnd
port 517 nsew
rlabel metal2 s 17658 18905 17766 19015 4 gnd
port 517 nsew
rlabel metal2 s 12186 22065 12294 22175 4 gnd
port 517 nsew
rlabel metal2 s 5946 2569 6054 2645 4 gnd
port 517 nsew
rlabel metal2 s 18426 19695 18534 19805 4 gnd
port 517 nsew
rlabel metal2 s 13914 1525 14022 1635 4 gnd
port 517 nsew
rlabel metal2 s 9690 1305 9798 1381 4 gnd
port 517 nsew
rlabel metal2 s 7674 13629 7782 13705 4 gnd
port 517 nsew
rlabel metal2 s 18426 12365 18534 12441 4 gnd
port 517 nsew
rlabel metal2 s 8442 6265 8550 6375 4 gnd
port 517 nsew
rlabel metal2 s 14682 7845 14790 7955 4 gnd
port 517 nsew
rlabel metal2 s 12186 25225 12294 25335 4 gnd
port 517 nsew
rlabel metal2 s 17658 16315 17766 16391 4 gnd
port 517 nsew
rlabel metal2 s 18426 23425 18534 23501 4 gnd
port 517 nsew
rlabel metal2 s 2682 1525 2790 1635 4 gnd
port 517 nsew
rlabel metal2 s 16410 15999 16518 16075 4 gnd
port 517 nsew
rlabel metal2 s 4698 3895 4806 4005 4 gnd
port 517 nsew
rlabel metal2 s 12666 21275 12774 21385 4 gnd
port 517 nsew
rlabel metal2 s 17178 19475 17286 19551 4 gnd
port 517 nsew
rlabel metal2 s 7674 17895 7782 17971 4 gnd
port 517 nsew
rlabel metal2 s 12666 3675 12774 3751 4 gnd
port 517 nsew
rlabel metal2 s 5178 20739 5286 20815 4 gnd
port 517 nsew
rlabel metal2 s 3450 13945 3558 14021 4 gnd
port 517 nsew
rlabel metal2 s 8442 18685 8550 18761 4 gnd
port 517 nsew
rlabel metal2 s 186 20265 294 20341 4 gnd
port 517 nsew
rlabel metal2 s 7674 5729 7782 5805 4 gnd
port 517 nsew
rlabel metal2 s 954 12365 1062 12441 4 gnd
port 517 nsew
rlabel metal2 s 5946 8889 6054 8965 4 gnd
port 517 nsew
rlabel metal2 s 9690 18685 9798 18761 4 gnd
port 517 nsew
rlabel metal2 s 10170 22065 10278 22175 4 gnd
port 517 nsew
rlabel metal2 s 8922 20739 9030 20815 4 gnd
port 517 nsew
rlabel metal2 s 11418 17895 11526 17971 4 gnd
port 517 nsew
rlabel metal2 s 12666 17579 12774 17655 4 gnd
port 517 nsew
rlabel metal2 s 954 8635 1062 8745 4 gnd
port 517 nsew
rlabel metal2 s 10938 8415 11046 8491 4 gnd
port 517 nsew
rlabel metal2 s 18906 12585 19014 12695 4 gnd
port 517 nsew
rlabel metal2 s 19674 23109 19782 23185 4 gnd
port 517 nsew
rlabel metal2 s 7674 16535 7782 16645 4 gnd
port 517 nsew
rlabel metal2 s 8922 10469 9030 10545 4 gnd
port 517 nsew
rlabel metal2 s 5946 21845 6054 21921 4 gnd
port 517 nsew
rlabel metal2 s 7674 17105 7782 17181 4 gnd
port 517 nsew
rlabel metal2 s 3450 7055 3558 7165 4 gnd
port 517 nsew
rlabel metal2 s 12666 20265 12774 20341 4 gnd
port 517 nsew
rlabel metal2 s 8442 23899 8550 23975 4 gnd
port 517 nsew
rlabel metal2 s 8922 19159 9030 19235 4 gnd
port 517 nsew
rlabel metal2 s 6426 2095 6534 2171 4 gnd
port 517 nsew
rlabel metal2 s 12186 7625 12294 7701 4 gnd
port 517 nsew
rlabel metal2 s 17178 24689 17286 24765 4 gnd
port 517 nsew
rlabel metal2 s 8922 5475 9030 5585 4 gnd
port 517 nsew
rlabel metal2 s 16410 9995 16518 10071 4 gnd
port 517 nsew
rlabel metal2 s 13914 23109 14022 23185 4 gnd
port 517 nsew
rlabel metal2 s 17178 11259 17286 11335 4 gnd
port 517 nsew
rlabel metal2 s 5178 3895 5286 4005 4 gnd
port 517 nsew
rlabel metal2 s 15162 13629 15270 13705 4 gnd
port 517 nsew
rlabel metal2 s 8922 13945 9030 14021 4 gnd
port 517 nsew
rlabel metal2 s 13434 4685 13542 4795 4 gnd
port 517 nsew
rlabel metal2 s 15162 5729 15270 5805 4 gnd
port 517 nsew
rlabel metal2 s 6426 735 6534 845 4 gnd
port 517 nsew
rlabel metal2 s 4698 11005 4806 11115 4 gnd
port 517 nsew
rlabel metal2 s 9690 515 9798 591 4 gnd
port 517 nsew
rlabel metal2 s 16410 6835 16518 6911 4 gnd
port 517 nsew
rlabel metal2 s 17658 12049 17766 12125 4 gnd
port 517 nsew
rlabel metal2 s 3450 16789 3558 16865 4 gnd
port 517 nsew
rlabel metal2 s 12186 11575 12294 11651 4 gnd
port 517 nsew
rlabel metal2 s 2682 3359 2790 3435 4 gnd
port 517 nsew
rlabel metal2 s 13914 17579 14022 17655 4 gnd
port 517 nsew
rlabel metal2 s 18906 14165 19014 14275 4 gnd
port 517 nsew
rlabel metal2 s 5946 25225 6054 25335 4 gnd
port 517 nsew
rlabel metal2 s 15930 21275 16038 21385 4 gnd
port 517 nsew
rlabel metal2 s 1434 3359 1542 3435 4 gnd
port 517 nsew
rlabel metal2 s 5178 1525 5286 1635 4 gnd
port 517 nsew
rlabel metal2 s 186 20739 294 20815 4 gnd
port 517 nsew
rlabel metal2 s 8922 3895 9030 4005 4 gnd
port 517 nsew
rlabel metal2 s 8442 20265 8550 20341 4 gnd
port 517 nsew
rlabel metal2 s 12666 17895 12774 17971 4 gnd
port 517 nsew
rlabel metal2 s 4698 14735 4806 14811 4 gnd
port 517 nsew
rlabel metal2 s 14682 16535 14790 16645 4 gnd
port 517 nsew
rlabel metal2 s 2202 23645 2310 23755 4 gnd
port 517 nsew
rlabel metal2 s 10170 2885 10278 2961 4 gnd
port 517 nsew
rlabel metal2 s 12666 13945 12774 14021 4 gnd
port 517 nsew
rlabel metal2 s 15930 20265 16038 20341 4 gnd
port 517 nsew
rlabel metal2 s 5178 19475 5286 19551 4 gnd
port 517 nsew
rlabel metal2 s 8442 16535 8550 16645 4 gnd
port 517 nsew
rlabel metal2 s 12186 22635 12294 22711 4 gnd
port 517 nsew
rlabel metal2 s 16410 13155 16518 13231 4 gnd
port 517 nsew
rlabel metal2 s 9690 15525 9798 15601 4 gnd
port 517 nsew
rlabel metal2 s 15162 11005 15270 11115 4 gnd
port 517 nsew
rlabel metal2 s 954 7055 1062 7165 4 gnd
port 517 nsew
rlabel metal2 s 4698 20265 4806 20341 4 gnd
port 517 nsew
rlabel metal2 s 5946 11005 6054 11115 4 gnd
port 517 nsew
rlabel metal2 s 18426 18115 18534 18225 4 gnd
port 517 nsew
rlabel metal2 s 17178 9995 17286 10071 4 gnd
port 517 nsew
rlabel metal2 s 18426 14419 18534 14495 4 gnd
port 517 nsew
rlabel metal2 s 12186 14165 12294 14275 4 gnd
port 517 nsew
rlabel metal2 s 14682 15999 14790 16075 4 gnd
port 517 nsew
rlabel metal2 s 3930 21845 4038 21921 4 gnd
port 517 nsew
rlabel metal2 s 3930 11795 4038 11905 4 gnd
port 517 nsew
rlabel metal2 s 10938 10469 11046 10545 4 gnd
port 517 nsew
rlabel metal2 s 5178 25225 5286 25335 4 gnd
port 517 nsew
rlabel metal2 s 12186 20265 12294 20341 4 gnd
port 517 nsew
rlabel metal2 s 3930 12049 4038 12125 4 gnd
port 517 nsew
rlabel metal2 s 13434 989 13542 1065 4 gnd
port 517 nsew
rlabel metal2 s 15930 3675 16038 3751 4 gnd
port 517 nsew
rlabel metal2 s 5946 4465 6054 4541 4 gnd
port 517 nsew
rlabel metal2 s 13914 23645 14022 23755 4 gnd
port 517 nsew
rlabel metal2 s 14682 18685 14790 18761 4 gnd
port 517 nsew
rlabel metal2 s 14682 25225 14790 25335 4 gnd
port 517 nsew
rlabel metal2 s 14682 7309 14790 7385 4 gnd
port 517 nsew
rlabel metal2 s 2682 4685 2790 4795 4 gnd
port 517 nsew
rlabel metal2 s 4698 3675 4806 3751 4 gnd
port 517 nsew
rlabel metal2 s 18426 10785 18534 10861 4 gnd
port 517 nsew
rlabel metal2 s 2682 6835 2790 6911 4 gnd
port 517 nsew
rlabel metal2 s 15930 25005 16038 25081 4 gnd
port 517 nsew
rlabel metal2 s 2202 18905 2310 19015 4 gnd
port 517 nsew
rlabel metal2 s 16410 16535 16518 16645 4 gnd
port 517 nsew
rlabel metal2 s 12186 2569 12294 2645 4 gnd
port 517 nsew
rlabel metal2 s 11418 20485 11526 20595 4 gnd
port 517 nsew
rlabel metal2 s 15162 12585 15270 12695 4 gnd
port 517 nsew
rlabel metal2 s 7674 22319 7782 22395 4 gnd
port 517 nsew
rlabel metal2 s 19674 18685 19782 18761 4 gnd
port 517 nsew
rlabel metal2 s 17658 989 17766 1065 4 gnd
port 517 nsew
rlabel metal2 s 4698 9679 4806 9755 4 gnd
port 517 nsew
rlabel metal2 s 6426 23425 6534 23501 4 gnd
port 517 nsew
rlabel metal2 s 14682 1525 14790 1635 4 gnd
port 517 nsew
rlabel metal2 s 954 14165 1062 14275 4 gnd
port 517 nsew
rlabel metal2 s 15162 7625 15270 7701 4 gnd
port 517 nsew
rlabel metal2 s 5946 20485 6054 20595 4 gnd
port 517 nsew
rlabel metal2 s 5946 23645 6054 23755 4 gnd
port 517 nsew
rlabel metal2 s 14682 8099 14790 8175 4 gnd
port 517 nsew
rlabel metal2 s 14682 16789 14790 16865 4 gnd
port 517 nsew
rlabel metal2 s 17658 14165 17766 14275 4 gnd
port 517 nsew
rlabel metal2 s 17178 9679 17286 9755 4 gnd
port 517 nsew
rlabel metal2 s 17178 13945 17286 14021 4 gnd
port 517 nsew
rlabel metal2 s 15930 12839 16038 12915 4 gnd
port 517 nsew
rlabel metal2 s 3930 8099 4038 8175 4 gnd
port 517 nsew
rlabel metal2 s 12186 7309 12294 7385 4 gnd
port 517 nsew
rlabel metal2 s 2202 18115 2310 18225 4 gnd
port 517 nsew
rlabel metal2 s 10938 515 11046 591 4 gnd
port 517 nsew
rlabel metal2 s 2202 14419 2310 14495 4 gnd
port 517 nsew
rlabel metal2 s 16410 6265 16518 6375 4 gnd
port 517 nsew
rlabel metal2 s 13434 20485 13542 20595 4 gnd
port 517 nsew
rlabel metal2 s 14682 4685 14790 4795 4 gnd
port 517 nsew
rlabel metal2 s 17178 14735 17286 14811 4 gnd
port 517 nsew
rlabel metal2 s 3930 8889 4038 8965 4 gnd
port 517 nsew
rlabel metal2 s 7674 23899 7782 23975 4 gnd
port 517 nsew
rlabel metal2 s 14682 9425 14790 9535 4 gnd
port 517 nsew
rlabel metal2 s 17178 515 17286 591 4 gnd
port 517 nsew
rlabel metal2 s 7194 23899 7302 23975 4 gnd
port 517 nsew
rlabel metal2 s 12186 21529 12294 21605 4 gnd
port 517 nsew
rlabel metal2 s 15162 515 15270 591 4 gnd
port 517 nsew
rlabel metal2 s 17658 6519 17766 6595 4 gnd
port 517 nsew
rlabel metal2 s 2682 21845 2790 21921 4 gnd
port 517 nsew
rlabel metal2 s 4698 9995 4806 10071 4 gnd
port 517 nsew
rlabel metal2 s 18426 989 18534 1065 4 gnd
port 517 nsew
rlabel metal2 s 12666 10469 12774 10545 4 gnd
port 517 nsew
rlabel metal2 s 8442 22319 8550 22395 4 gnd
port 517 nsew
rlabel metal2 s 13914 2569 14022 2645 4 gnd
port 517 nsew
rlabel metal2 s 3930 16789 4038 16865 4 gnd
port 517 nsew
rlabel metal2 s 5946 1525 6054 1635 4 gnd
port 517 nsew
rlabel metal2 s 15162 2315 15270 2425 4 gnd
port 517 nsew
rlabel metal2 s 14682 11575 14790 11651 4 gnd
port 517 nsew
rlabel metal2 s 186 199 294 275 4 gnd
port 517 nsew
rlabel metal2 s 13434 14955 13542 15065 4 gnd
port 517 nsew
rlabel metal2 s 5178 23645 5286 23755 4 gnd
port 517 nsew
rlabel metal2 s 15162 1525 15270 1635 4 gnd
port 517 nsew
rlabel metal2 s 5946 7845 6054 7955 4 gnd
port 517 nsew
rlabel metal2 s 7194 25225 7302 25335 4 gnd
port 517 nsew
rlabel metal2 s 9690 10469 9798 10545 4 gnd
port 517 nsew
rlabel metal2 s 10938 19475 11046 19551 4 gnd
port 517 nsew
rlabel metal2 s 19674 1779 19782 1855 4 gnd
port 517 nsew
rlabel metal2 s 954 9995 1062 10071 4 gnd
port 517 nsew
rlabel metal2 s 3930 12365 4038 12441 4 gnd
port 517 nsew
rlabel metal2 s 3930 21055 4038 21131 4 gnd
port 517 nsew
rlabel metal2 s 12666 8099 12774 8175 4 gnd
port 517 nsew
rlabel metal2 s 5946 17325 6054 17435 4 gnd
port 517 nsew
rlabel metal2 s 17178 21845 17286 21921 4 gnd
port 517 nsew
rlabel metal2 s 3930 989 4038 1065 4 gnd
port 517 nsew
rlabel metal2 s 7194 6045 7302 6121 4 gnd
port 517 nsew
rlabel metal2 s 6426 17579 6534 17655 4 gnd
port 517 nsew
rlabel metal2 s 186 13945 294 14021 4 gnd
port 517 nsew
rlabel metal2 s 7674 13155 7782 13231 4 gnd
port 517 nsew
rlabel metal2 s 16410 10785 16518 10861 4 gnd
port 517 nsew
rlabel metal2 s 13434 13375 13542 13485 4 gnd
port 517 nsew
rlabel metal2 s 12666 23425 12774 23501 4 gnd
port 517 nsew
rlabel metal2 s 11418 21055 11526 21131 4 gnd
port 517 nsew
rlabel metal2 s 14682 21055 14790 21131 4 gnd
port 517 nsew
rlabel metal2 s 10170 14165 10278 14275 4 gnd
port 517 nsew
rlabel metal2 s 18906 19475 19014 19551 4 gnd
port 517 nsew
rlabel metal2 s 13914 14955 14022 15065 4 gnd
port 517 nsew
rlabel metal2 s 14682 11795 14790 11905 4 gnd
port 517 nsew
rlabel metal2 s 11418 23109 11526 23185 4 gnd
port 517 nsew
rlabel metal2 s 2202 6835 2310 6911 4 gnd
port 517 nsew
rlabel metal2 s 14682 14419 14790 14495 4 gnd
port 517 nsew
rlabel metal2 s 186 6265 294 6375 4 gnd
port 517 nsew
rlabel metal2 s 5178 18369 5286 18445 4 gnd
port 517 nsew
rlabel metal2 s 9690 2095 9798 2171 4 gnd
port 517 nsew
rlabel metal2 s 11418 8415 11526 8491 4 gnd
port 517 nsew
rlabel metal2 s 954 18115 1062 18225 4 gnd
port 517 nsew
rlabel metal2 s 12666 24215 12774 24291 4 gnd
port 517 nsew
rlabel metal2 s 18426 19159 18534 19235 4 gnd
port 517 nsew
rlabel metal2 s 2202 10785 2310 10861 4 gnd
port 517 nsew
rlabel metal2 s 186 21529 294 21605 4 gnd
port 517 nsew
rlabel metal2 s 4698 19695 4806 19805 4 gnd
port 517 nsew
rlabel metal2 s 11418 16789 11526 16865 4 gnd
port 517 nsew
rlabel metal2 s 18906 12839 19014 12915 4 gnd
port 517 nsew
rlabel metal2 s 8442 13155 8550 13231 4 gnd
port 517 nsew
rlabel metal2 s 18426 22855 18534 22965 4 gnd
port 517 nsew
rlabel metal2 s 186 6519 294 6595 4 gnd
port 517 nsew
rlabel metal2 s 2202 7309 2310 7385 4 gnd
port 517 nsew
rlabel metal2 s 1434 8415 1542 8491 4 gnd
port 517 nsew
rlabel metal2 s 2682 735 2790 845 4 gnd
port 517 nsew
rlabel metal2 s 13434 25005 13542 25081 4 gnd
port 517 nsew
rlabel metal2 s 6426 13375 6534 13485 4 gnd
port 517 nsew
rlabel metal2 s 6426 11259 6534 11335 4 gnd
port 517 nsew
rlabel metal2 s 15162 14955 15270 15065 4 gnd
port 517 nsew
rlabel metal2 s 18906 735 19014 845 4 gnd
port 517 nsew
rlabel metal2 s 8922 4149 9030 4225 4 gnd
port 517 nsew
rlabel metal2 s 15162 15209 15270 15285 4 gnd
port 517 nsew
rlabel metal2 s 6426 14419 6534 14495 4 gnd
port 517 nsew
rlabel metal2 s 9690 12839 9798 12915 4 gnd
port 517 nsew
rlabel metal2 s 186 3105 294 3215 4 gnd
port 517 nsew
rlabel metal2 s 4698 24689 4806 24765 4 gnd
port 517 nsew
rlabel metal2 s 13914 9679 14022 9755 4 gnd
port 517 nsew
rlabel metal2 s 7674 13375 7782 13485 4 gnd
port 517 nsew
rlabel metal2 s 8442 16789 8550 16865 4 gnd
port 517 nsew
rlabel metal2 s 2682 13375 2790 13485 4 gnd
port 517 nsew
rlabel metal2 s 19674 18115 19782 18225 4 gnd
port 517 nsew
rlabel metal2 s 16410 3105 16518 3215 4 gnd
port 517 nsew
rlabel metal2 s 13914 10785 14022 10861 4 gnd
port 517 nsew
rlabel metal2 s 2202 15209 2310 15285 4 gnd
port 517 nsew
rlabel metal2 s 17178 10785 17286 10861 4 gnd
port 517 nsew
rlabel metal2 s 18906 6265 19014 6375 4 gnd
port 517 nsew
rlabel metal2 s 8922 199 9030 275 4 gnd
port 517 nsew
rlabel metal2 s 16410 9425 16518 9535 4 gnd
port 517 nsew
rlabel metal2 s 9690 19159 9798 19235 4 gnd
port 517 nsew
rlabel metal2 s 11418 8889 11526 8965 4 gnd
port 517 nsew
rlabel metal2 s 2682 23109 2790 23185 4 gnd
port 517 nsew
rlabel metal2 s 5178 14165 5286 14275 4 gnd
port 517 nsew
rlabel metal2 s 186 1525 294 1635 4 gnd
port 517 nsew
rlabel metal2 s 18906 8635 19014 8745 4 gnd
port 517 nsew
rlabel metal2 s 14682 17105 14790 17181 4 gnd
port 517 nsew
rlabel metal2 s 15930 14165 16038 14275 4 gnd
port 517 nsew
rlabel metal2 s 5178 6519 5286 6595 4 gnd
port 517 nsew
rlabel metal2 s 14682 6835 14790 6911 4 gnd
port 517 nsew
rlabel metal2 s 5178 1305 5286 1381 4 gnd
port 517 nsew
rlabel metal2 s 8442 1305 8550 1381 4 gnd
port 517 nsew
rlabel metal2 s 10170 515 10278 591 4 gnd
port 517 nsew
rlabel metal2 s 1434 18115 1542 18225 4 gnd
port 517 nsew
rlabel metal2 s 9690 3895 9798 4005 4 gnd
port 517 nsew
rlabel metal2 s 6426 11575 6534 11651 4 gnd
port 517 nsew
rlabel metal2 s 9690 21529 9798 21605 4 gnd
port 517 nsew
rlabel metal2 s 19674 8635 19782 8745 4 gnd
port 517 nsew
rlabel metal2 s 15930 8635 16038 8745 4 gnd
port 517 nsew
rlabel metal2 s 2202 8889 2310 8965 4 gnd
port 517 nsew
rlabel metal2 s 2682 24435 2790 24545 4 gnd
port 517 nsew
rlabel metal2 s 10938 11575 11046 11651 4 gnd
port 517 nsew
rlabel metal2 s 16410 25225 16518 25335 4 gnd
port 517 nsew
rlabel metal2 s 3450 5729 3558 5805 4 gnd
port 517 nsew
rlabel metal2 s 6426 1525 6534 1635 4 gnd
port 517 nsew
rlabel metal2 s 1434 21529 1542 21605 4 gnd
port 517 nsew
rlabel metal2 s 13434 15745 13542 15855 4 gnd
port 517 nsew
rlabel metal2 s 19674 8099 19782 8175 4 gnd
port 517 nsew
rlabel metal2 s 8442 3675 8550 3751 4 gnd
port 517 nsew
rlabel metal2 s 12186 5255 12294 5331 4 gnd
port 517 nsew
rlabel metal2 s 19674 13375 19782 13485 4 gnd
port 517 nsew
rlabel metal2 s 18906 9425 19014 9535 4 gnd
port 517 nsew
rlabel metal2 s 1434 1525 1542 1635 4 gnd
port 517 nsew
rlabel metal2 s 17178 16535 17286 16645 4 gnd
port 517 nsew
rlabel metal2 s 8922 9995 9030 10071 4 gnd
port 517 nsew
rlabel metal2 s 7194 10215 7302 10325 4 gnd
port 517 nsew
rlabel metal2 s 7674 22635 7782 22711 4 gnd
port 517 nsew
rlabel metal2 s 186 14419 294 14495 4 gnd
port 517 nsew
rlabel metal2 s 18906 23109 19014 23185 4 gnd
port 517 nsew
rlabel metal2 s 8442 14419 8550 14495 4 gnd
port 517 nsew
rlabel metal2 s 13434 5729 13542 5805 4 gnd
port 517 nsew
rlabel metal2 s 12186 19949 12294 20025 4 gnd
port 517 nsew
rlabel metal2 s 16410 23645 16518 23755 4 gnd
port 517 nsew
rlabel metal2 s 3930 15745 4038 15855 4 gnd
port 517 nsew
rlabel metal2 s 4698 15209 4806 15285 4 gnd
port 517 nsew
rlabel metal2 s 9690 19695 9798 19805 4 gnd
port 517 nsew
rlabel metal2 s 13914 7309 14022 7385 4 gnd
port 517 nsew
rlabel metal2 s 7674 15209 7782 15285 4 gnd
port 517 nsew
rlabel metal2 s 3450 18685 3558 18761 4 gnd
port 517 nsew
rlabel metal2 s 8442 17325 8550 17435 4 gnd
port 517 nsew
rlabel metal2 s 3930 16315 4038 16391 4 gnd
port 517 nsew
rlabel metal2 s 10938 3895 11046 4005 4 gnd
port 517 nsew
rlabel metal2 s 3930 17325 4038 17435 4 gnd
port 517 nsew
rlabel metal2 s 8922 3359 9030 3435 4 gnd
port 517 nsew
rlabel metal2 s 15930 4939 16038 5015 4 gnd
port 517 nsew
rlabel metal2 s 1434 8889 1542 8965 4 gnd
port 517 nsew
rlabel metal2 s 3450 8415 3558 8491 4 gnd
port 517 nsew
rlabel metal2 s 2202 11575 2310 11651 4 gnd
port 517 nsew
rlabel metal2 s 6426 8099 6534 8175 4 gnd
port 517 nsew
rlabel metal2 s 12666 1525 12774 1635 4 gnd
port 517 nsew
rlabel metal2 s 2202 11795 2310 11905 4 gnd
port 517 nsew
rlabel metal2 s 17658 12839 17766 12915 4 gnd
port 517 nsew
rlabel metal2 s 7194 14165 7302 14275 4 gnd
port 517 nsew
rlabel metal2 s 10938 18685 11046 18761 4 gnd
port 517 nsew
rlabel metal2 s 10938 199 11046 275 4 gnd
port 517 nsew
rlabel metal2 s 10938 20265 11046 20341 4 gnd
port 517 nsew
rlabel metal2 s 17178 14419 17286 14495 4 gnd
port 517 nsew
rlabel metal2 s 5946 23899 6054 23975 4 gnd
port 517 nsew
rlabel metal2 s 10938 5729 11046 5805 4 gnd
port 517 nsew
rlabel metal2 s 4698 19475 4806 19551 4 gnd
port 517 nsew
rlabel metal2 s 17178 2095 17286 2171 4 gnd
port 517 nsew
rlabel metal2 s 15930 12585 16038 12695 4 gnd
port 517 nsew
rlabel metal2 s 3930 17579 4038 17655 4 gnd
port 517 nsew
rlabel metal2 s 9690 6265 9798 6375 4 gnd
port 517 nsew
rlabel metal2 s 7674 735 7782 845 4 gnd
port 517 nsew
rlabel metal2 s 16410 16315 16518 16391 4 gnd
port 517 nsew
rlabel metal2 s 12666 11575 12774 11651 4 gnd
port 517 nsew
rlabel metal2 s 3450 7309 3558 7385 4 gnd
port 517 nsew
rlabel metal2 s 7194 14735 7302 14811 4 gnd
port 517 nsew
rlabel metal2 s 3450 6265 3558 6375 4 gnd
port 517 nsew
rlabel metal2 s 954 17325 1062 17435 4 gnd
port 517 nsew
rlabel metal2 s 17658 6045 17766 6121 4 gnd
port 517 nsew
rlabel metal2 s 18426 20485 18534 20595 4 gnd
port 517 nsew
rlabel metal2 s 18906 9205 19014 9281 4 gnd
port 517 nsew
rlabel metal2 s 7194 11575 7302 11651 4 gnd
port 517 nsew
rlabel metal2 s 17658 9425 17766 9535 4 gnd
port 517 nsew
rlabel metal2 s 3450 24689 3558 24765 4 gnd
port 517 nsew
rlabel metal2 s 17178 989 17286 1065 4 gnd
port 517 nsew
rlabel metal2 s 17658 25225 17766 25335 4 gnd
port 517 nsew
rlabel metal2 s 16410 18685 16518 18761 4 gnd
port 517 nsew
rlabel metal2 s 2202 6519 2310 6595 4 gnd
port 517 nsew
rlabel metal2 s 17658 4149 17766 4225 4 gnd
port 517 nsew
rlabel metal2 s 15930 11795 16038 11905 4 gnd
port 517 nsew
rlabel metal2 s 10938 2315 11046 2425 4 gnd
port 517 nsew
rlabel metal2 s 11418 20265 11526 20341 4 gnd
port 517 nsew
rlabel metal2 s 8922 15999 9030 16075 4 gnd
port 517 nsew
rlabel metal2 s 17658 16535 17766 16645 4 gnd
port 517 nsew
rlabel metal2 s 10170 2095 10278 2171 4 gnd
port 517 nsew
rlabel metal2 s 10170 12049 10278 12125 4 gnd
port 517 nsew
rlabel metal2 s 18426 9679 18534 9755 4 gnd
port 517 nsew
rlabel metal2 s 6426 6835 6534 6911 4 gnd
port 517 nsew
rlabel metal2 s 954 20485 1062 20595 4 gnd
port 517 nsew
rlabel metal2 s 7194 3895 7302 4005 4 gnd
port 517 nsew
rlabel metal2 s 2682 22855 2790 22965 4 gnd
port 517 nsew
rlabel metal2 s 186 21275 294 21385 4 gnd
port 517 nsew
rlabel metal2 s 186 2315 294 2425 4 gnd
port 517 nsew
rlabel metal2 s 15162 2569 15270 2645 4 gnd
port 517 nsew
rlabel metal2 s 15930 3895 16038 4005 4 gnd
port 517 nsew
rlabel metal2 s 14682 21529 14790 21605 4 gnd
port 517 nsew
rlabel metal2 s 3450 23109 3558 23185 4 gnd
port 517 nsew
rlabel metal2 s 7674 20265 7782 20341 4 gnd
port 517 nsew
rlabel metal2 s 12666 25225 12774 25335 4 gnd
port 517 nsew
rlabel metal2 s 12186 23899 12294 23975 4 gnd
port 517 nsew
rlabel metal2 s 13434 735 13542 845 4 gnd
port 517 nsew
rlabel metal2 s 5178 12839 5286 12915 4 gnd
port 517 nsew
rlabel metal2 s 13434 25225 13542 25335 4 gnd
port 517 nsew
rlabel metal2 s 15162 14165 15270 14275 4 gnd
port 517 nsew
rlabel metal2 s 10170 17325 10278 17435 4 gnd
port 517 nsew
rlabel metal2 s 16410 11005 16518 11115 4 gnd
port 517 nsew
rlabel metal2 s 19674 17325 19782 17435 4 gnd
port 517 nsew
rlabel metal2 s 10938 17105 11046 17181 4 gnd
port 517 nsew
rlabel metal2 s 13914 18369 14022 18445 4 gnd
port 517 nsew
rlabel metal2 s 2682 9995 2790 10071 4 gnd
port 517 nsew
rlabel metal2 s 5178 7625 5286 7701 4 gnd
port 517 nsew
rlabel metal2 s 12186 15209 12294 15285 4 gnd
port 517 nsew
rlabel metal2 s 4698 20739 4806 20815 4 gnd
port 517 nsew
rlabel metal2 s 15930 5475 16038 5585 4 gnd
port 517 nsew
rlabel metal2 s 9690 4685 9798 4795 4 gnd
port 517 nsew
rlabel metal2 s 13914 12585 14022 12695 4 gnd
port 517 nsew
rlabel metal2 s 18906 14735 19014 14811 4 gnd
port 517 nsew
rlabel metal2 s 18426 7625 18534 7701 4 gnd
port 517 nsew
rlabel metal2 s 954 10785 1062 10861 4 gnd
port 517 nsew
rlabel metal2 s 6426 22319 6534 22395 4 gnd
port 517 nsew
rlabel metal2 s 10938 9205 11046 9281 4 gnd
port 517 nsew
rlabel metal2 s 7194 13375 7302 13485 4 gnd
port 517 nsew
rlabel metal2 s 186 17325 294 17435 4 gnd
port 517 nsew
rlabel metal2 s 19674 6519 19782 6595 4 gnd
port 517 nsew
rlabel metal2 s 10170 19475 10278 19551 4 gnd
port 517 nsew
rlabel metal2 s 3450 19475 3558 19551 4 gnd
port 517 nsew
rlabel metal2 s 12666 6835 12774 6911 4 gnd
port 517 nsew
rlabel metal2 s 13914 18115 14022 18225 4 gnd
port 517 nsew
rlabel metal2 s 2202 23899 2310 23975 4 gnd
port 517 nsew
rlabel metal2 s 3450 4149 3558 4225 4 gnd
port 517 nsew
rlabel metal2 s 2682 16315 2790 16391 4 gnd
port 517 nsew
rlabel metal2 s 3930 4685 4038 4795 4 gnd
port 517 nsew
rlabel metal2 s 18906 7309 19014 7385 4 gnd
port 517 nsew
rlabel metal2 s 15930 8415 16038 8491 4 gnd
port 517 nsew
rlabel metal2 s 5178 20265 5286 20341 4 gnd
port 517 nsew
rlabel metal2 s 7674 12365 7782 12441 4 gnd
port 517 nsew
rlabel metal2 s 18906 13945 19014 14021 4 gnd
port 517 nsew
rlabel metal2 s 15162 24689 15270 24765 4 gnd
port 517 nsew
rlabel metal2 s 10938 7309 11046 7385 4 gnd
port 517 nsew
rlabel metal2 s 10938 21529 11046 21605 4 gnd
port 517 nsew
rlabel metal2 s 11418 2315 11526 2425 4 gnd
port 517 nsew
rlabel metal2 s 15930 14419 16038 14495 4 gnd
port 517 nsew
rlabel metal2 s 11418 13375 11526 13485 4 gnd
port 517 nsew
rlabel metal2 s 1434 15209 1542 15285 4 gnd
port 517 nsew
rlabel metal2 s 8442 14165 8550 14275 4 gnd
port 517 nsew
rlabel metal2 s 9690 15745 9798 15855 4 gnd
port 517 nsew
rlabel metal2 s 5946 23425 6054 23501 4 gnd
port 517 nsew
rlabel metal2 s 15930 13945 16038 14021 4 gnd
port 517 nsew
rlabel metal2 s 2202 14165 2310 14275 4 gnd
port 517 nsew
rlabel metal2 s 8442 13629 8550 13705 4 gnd
port 517 nsew
rlabel metal2 s 186 19949 294 20025 4 gnd
port 517 nsew
rlabel metal2 s 13914 5729 14022 5805 4 gnd
port 517 nsew
rlabel metal2 s 16410 15209 16518 15285 4 gnd
port 517 nsew
rlabel metal2 s 17658 5255 17766 5331 4 gnd
port 517 nsew
rlabel metal2 s 13434 18685 13542 18761 4 gnd
port 517 nsew
rlabel metal2 s 5946 11575 6054 11651 4 gnd
port 517 nsew
rlabel metal2 s 15930 15999 16038 16075 4 gnd
port 517 nsew
rlabel metal2 s 2682 7625 2790 7701 4 gnd
port 517 nsew
rlabel metal2 s 17658 15209 17766 15285 4 gnd
port 517 nsew
rlabel metal2 s 3930 14955 4038 15065 4 gnd
port 517 nsew
rlabel metal2 s 12186 13629 12294 13705 4 gnd
port 517 nsew
rlabel metal2 s 2682 11795 2790 11905 4 gnd
port 517 nsew
rlabel metal2 s 2682 23645 2790 23755 4 gnd
port 517 nsew
rlabel metal2 s 6426 515 6534 591 4 gnd
port 517 nsew
rlabel metal2 s 10938 5255 11046 5331 4 gnd
port 517 nsew
rlabel metal2 s 5178 20485 5286 20595 4 gnd
port 517 nsew
rlabel metal2 s 14682 2569 14790 2645 4 gnd
port 517 nsew
rlabel metal2 s 4698 17579 4806 17655 4 gnd
port 517 nsew
rlabel metal2 s 4698 2885 4806 2961 4 gnd
port 517 nsew
rlabel metal2 s 6426 13945 6534 14021 4 gnd
port 517 nsew
rlabel metal2 s 6426 19159 6534 19235 4 gnd
port 517 nsew
rlabel metal2 s 4698 989 4806 1065 4 gnd
port 517 nsew
rlabel metal2 s 13914 17325 14022 17435 4 gnd
port 517 nsew
rlabel metal2 s 14682 13375 14790 13485 4 gnd
port 517 nsew
rlabel metal2 s 7194 5475 7302 5585 4 gnd
port 517 nsew
rlabel metal2 s 6426 22855 6534 22965 4 gnd
port 517 nsew
rlabel metal2 s 7674 2885 7782 2961 4 gnd
port 517 nsew
rlabel metal2 s 12186 10215 12294 10325 4 gnd
port 517 nsew
rlabel metal2 s 18906 5255 19014 5331 4 gnd
port 517 nsew
rlabel metal2 s 1434 16315 1542 16391 4 gnd
port 517 nsew
rlabel metal2 s 954 14955 1062 15065 4 gnd
port 517 nsew
rlabel metal2 s 18426 15999 18534 16075 4 gnd
port 517 nsew
rlabel metal2 s 12666 18685 12774 18761 4 gnd
port 517 nsew
rlabel metal2 s 954 -55 1062 55 4 gnd
port 517 nsew
rlabel metal2 s 13914 3895 14022 4005 4 gnd
port 517 nsew
rlabel metal2 s 954 3895 1062 4005 4 gnd
port 517 nsew
rlabel metal2 s 12186 8099 12294 8175 4 gnd
port 517 nsew
rlabel metal2 s 15930 24435 16038 24545 4 gnd
port 517 nsew
rlabel metal2 s 7194 23645 7302 23755 4 gnd
port 517 nsew
rlabel metal2 s 17658 23645 17766 23755 4 gnd
port 517 nsew
rlabel metal2 s 6426 23645 6534 23755 4 gnd
port 517 nsew
rlabel metal2 s 10938 4685 11046 4795 4 gnd
port 517 nsew
rlabel metal2 s 18426 24435 18534 24545 4 gnd
port 517 nsew
rlabel metal2 s 16410 22319 16518 22395 4 gnd
port 517 nsew
rlabel metal2 s 17658 3359 17766 3435 4 gnd
port 517 nsew
rlabel metal2 s 17658 7055 17766 7165 4 gnd
port 517 nsew
rlabel metal2 s 12186 8889 12294 8965 4 gnd
port 517 nsew
rlabel metal2 s 186 17105 294 17181 4 gnd
port 517 nsew
rlabel metal2 s 8442 17579 8550 17655 4 gnd
port 517 nsew
rlabel metal2 s 1434 735 1542 845 4 gnd
port 517 nsew
rlabel metal2 s 17658 22065 17766 22175 4 gnd
port 517 nsew
rlabel metal2 s 11418 11575 11526 11651 4 gnd
port 517 nsew
rlabel metal2 s 18426 2315 18534 2425 4 gnd
port 517 nsew
rlabel metal2 s 13914 17105 14022 17181 4 gnd
port 517 nsew
rlabel metal2 s 186 24689 294 24765 4 gnd
port 517 nsew
rlabel metal2 s 7194 20739 7302 20815 4 gnd
port 517 nsew
rlabel metal2 s 6426 19475 6534 19551 4 gnd
port 517 nsew
rlabel metal2 s 13434 22065 13542 22175 4 gnd
port 517 nsew
rlabel metal2 s 5946 9679 6054 9755 4 gnd
port 517 nsew
rlabel metal2 s 13434 14419 13542 14495 4 gnd
port 517 nsew
rlabel metal2 s 18426 515 18534 591 4 gnd
port 517 nsew
rlabel metal2 s 1434 19475 1542 19551 4 gnd
port 517 nsew
rlabel metal2 s 13434 17579 13542 17655 4 gnd
port 517 nsew
rlabel metal2 s 13434 1305 13542 1381 4 gnd
port 517 nsew
rlabel metal2 s 3450 23645 3558 23755 4 gnd
port 517 nsew
rlabel metal2 s 8922 6519 9030 6595 4 gnd
port 517 nsew
rlabel metal2 s 2682 14955 2790 15065 4 gnd
port 517 nsew
rlabel metal2 s 10170 8889 10278 8965 4 gnd
port 517 nsew
rlabel metal2 s 17178 16315 17286 16391 4 gnd
port 517 nsew
rlabel metal2 s 3450 13375 3558 13485 4 gnd
port 517 nsew
rlabel metal2 s 19674 6045 19782 6121 4 gnd
port 517 nsew
rlabel metal2 s 11418 15745 11526 15855 4 gnd
port 517 nsew
rlabel metal2 s 8922 14419 9030 14495 4 gnd
port 517 nsew
rlabel metal2 s 3930 10215 4038 10325 4 gnd
port 517 nsew
rlabel metal2 s 3450 10215 3558 10325 4 gnd
port 517 nsew
rlabel metal2 s 13914 989 14022 1065 4 gnd
port 517 nsew
rlabel metal2 s 14682 -55 14790 55 4 gnd
port 517 nsew
rlabel metal2 s 8442 21275 8550 21385 4 gnd
port 517 nsew
rlabel metal2 s 17658 19949 17766 20025 4 gnd
port 517 nsew
rlabel metal2 s 17658 3105 17766 3215 4 gnd
port 517 nsew
rlabel metal2 s 2682 15525 2790 15601 4 gnd
port 517 nsew
rlabel metal2 s 3930 2095 4038 2171 4 gnd
port 517 nsew
rlabel metal2 s 7674 21275 7782 21385 4 gnd
port 517 nsew
rlabel metal2 s 1434 4149 1542 4225 4 gnd
port 517 nsew
rlabel metal2 s 13434 10785 13542 10861 4 gnd
port 517 nsew
rlabel metal2 s 17178 3359 17286 3435 4 gnd
port 517 nsew
rlabel metal2 s 5946 12365 6054 12441 4 gnd
port 517 nsew
rlabel metal2 s 10170 25225 10278 25335 4 gnd
port 517 nsew
rlabel metal2 s 3930 3895 4038 4005 4 gnd
port 517 nsew
rlabel metal2 s 1434 21845 1542 21921 4 gnd
port 517 nsew
rlabel metal2 s 3450 14419 3558 14495 4 gnd
port 517 nsew
rlabel metal2 s 12666 7625 12774 7701 4 gnd
port 517 nsew
rlabel metal2 s 19674 20265 19782 20341 4 gnd
port 517 nsew
rlabel metal2 s 17658 15525 17766 15601 4 gnd
port 517 nsew
rlabel metal2 s 17178 15999 17286 16075 4 gnd
port 517 nsew
rlabel metal2 s 18426 3359 18534 3435 4 gnd
port 517 nsew
rlabel metal2 s 11418 9679 11526 9755 4 gnd
port 517 nsew
rlabel metal2 s 7674 11575 7782 11651 4 gnd
port 517 nsew
rlabel metal2 s 4698 23109 4806 23185 4 gnd
port 517 nsew
rlabel metal2 s 18906 5475 19014 5585 4 gnd
port 517 nsew
rlabel metal2 s 13434 7845 13542 7955 4 gnd
port 517 nsew
rlabel metal2 s 8922 21529 9030 21605 4 gnd
port 517 nsew
rlabel metal2 s 13434 17325 13542 17435 4 gnd
port 517 nsew
rlabel metal2 s 18426 20739 18534 20815 4 gnd
port 517 nsew
rlabel metal2 s 14682 21845 14790 21921 4 gnd
port 517 nsew
rlabel metal2 s 7194 23109 7302 23185 4 gnd
port 517 nsew
rlabel metal2 s 2202 3675 2310 3751 4 gnd
port 517 nsew
rlabel metal2 s 5178 9205 5286 9281 4 gnd
port 517 nsew
rlabel metal2 s 12186 2315 12294 2425 4 gnd
port 517 nsew
rlabel metal2 s 12666 735 12774 845 4 gnd
port 517 nsew
rlabel metal2 s 15162 9679 15270 9755 4 gnd
port 517 nsew
rlabel metal2 s 17658 22635 17766 22711 4 gnd
port 517 nsew
rlabel metal2 s 18426 10469 18534 10545 4 gnd
port 517 nsew
rlabel metal2 s 9690 6045 9798 6121 4 gnd
port 517 nsew
rlabel metal2 s 1434 6265 1542 6375 4 gnd
port 517 nsew
rlabel metal2 s 3450 16535 3558 16645 4 gnd
port 517 nsew
rlabel metal2 s 8922 12365 9030 12441 4 gnd
port 517 nsew
rlabel metal2 s 7194 19475 7302 19551 4 gnd
port 517 nsew
rlabel metal2 s 5178 14419 5286 14495 4 gnd
port 517 nsew
rlabel metal2 s 2202 3105 2310 3215 4 gnd
port 517 nsew
rlabel metal2 s 11418 14165 11526 14275 4 gnd
port 517 nsew
rlabel metal2 s 12666 22855 12774 22965 4 gnd
port 517 nsew
rlabel metal2 s 14682 5255 14790 5331 4 gnd
port 517 nsew
rlabel metal2 s 12666 15745 12774 15855 4 gnd
port 517 nsew
rlabel metal2 s 10170 6835 10278 6911 4 gnd
port 517 nsew
rlabel metal2 s 954 23425 1062 23501 4 gnd
port 517 nsew
rlabel metal2 s 10170 4465 10278 4541 4 gnd
port 517 nsew
rlabel metal2 s 10938 15999 11046 16075 4 gnd
port 517 nsew
rlabel metal2 s 1434 13629 1542 13705 4 gnd
port 517 nsew
rlabel metal2 s 17178 15745 17286 15855 4 gnd
port 517 nsew
rlabel metal2 s 7674 1525 7782 1635 4 gnd
port 517 nsew
rlabel metal2 s 1434 21055 1542 21131 4 gnd
port 517 nsew
rlabel metal2 s 5946 8415 6054 8491 4 gnd
port 517 nsew
rlabel metal2 s 17178 2569 17286 2645 4 gnd
port 517 nsew
rlabel metal2 s 16410 17105 16518 17181 4 gnd
port 517 nsew
rlabel metal2 s 15930 22855 16038 22965 4 gnd
port 517 nsew
rlabel metal2 s 3450 14955 3558 15065 4 gnd
port 517 nsew
rlabel metal2 s 9690 10785 9798 10861 4 gnd
port 517 nsew
rlabel metal2 s 13914 16535 14022 16645 4 gnd
port 517 nsew
rlabel metal2 s 3930 6519 4038 6595 4 gnd
port 517 nsew
rlabel metal2 s 19674 6835 19782 6911 4 gnd
port 517 nsew
rlabel metal2 s 10170 1305 10278 1381 4 gnd
port 517 nsew
rlabel metal2 s 13914 19949 14022 20025 4 gnd
port 517 nsew
rlabel metal2 s 186 23425 294 23501 4 gnd
port 517 nsew
rlabel metal2 s 5178 5255 5286 5331 4 gnd
port 517 nsew
rlabel metal2 s 3930 22855 4038 22965 4 gnd
port 517 nsew
rlabel metal2 s 186 11259 294 11335 4 gnd
port 517 nsew
rlabel metal2 s 15930 17105 16038 17181 4 gnd
port 517 nsew
rlabel metal2 s 17178 22855 17286 22965 4 gnd
port 517 nsew
rlabel metal2 s 13914 20485 14022 20595 4 gnd
port 517 nsew
rlabel metal2 s 2682 2095 2790 2171 4 gnd
port 517 nsew
rlabel metal2 s 17178 13155 17286 13231 4 gnd
port 517 nsew
rlabel metal2 s 18426 3105 18534 3215 4 gnd
port 517 nsew
rlabel metal2 s 2682 22635 2790 22711 4 gnd
port 517 nsew
rlabel metal2 s 10938 22855 11046 22965 4 gnd
port 517 nsew
rlabel metal2 s 6426 21845 6534 21921 4 gnd
port 517 nsew
rlabel metal2 s 8442 2569 8550 2645 4 gnd
port 517 nsew
rlabel metal2 s 12186 9679 12294 9755 4 gnd
port 517 nsew
rlabel metal2 s 186 5255 294 5331 4 gnd
port 517 nsew
rlabel metal2 s 8442 19159 8550 19235 4 gnd
port 517 nsew
rlabel metal2 s 18426 19475 18534 19551 4 gnd
port 517 nsew
rlabel metal2 s 10938 3675 11046 3751 4 gnd
port 517 nsew
rlabel metal2 s 14682 24689 14790 24765 4 gnd
port 517 nsew
rlabel metal2 s 19674 11005 19782 11115 4 gnd
port 517 nsew
rlabel metal2 s 9690 19949 9798 20025 4 gnd
port 517 nsew
rlabel metal2 s 6426 16315 6534 16391 4 gnd
port 517 nsew
rlabel metal2 s 17178 17325 17286 17435 4 gnd
port 517 nsew
rlabel metal2 s 3930 11005 4038 11115 4 gnd
port 517 nsew
rlabel metal2 s 3450 22635 3558 22711 4 gnd
port 517 nsew
rlabel metal2 s 3930 1525 4038 1635 4 gnd
port 517 nsew
rlabel metal2 s 17178 21275 17286 21385 4 gnd
port 517 nsew
rlabel metal2 s 18906 3359 19014 3435 4 gnd
port 517 nsew
rlabel metal2 s 7194 7625 7302 7701 4 gnd
port 517 nsew
rlabel metal2 s 9690 17895 9798 17971 4 gnd
port 517 nsew
rlabel metal2 s 11418 24215 11526 24291 4 gnd
port 517 nsew
rlabel metal2 s 9690 12585 9798 12695 4 gnd
port 517 nsew
rlabel metal2 s 10938 6265 11046 6375 4 gnd
port 517 nsew
rlabel metal2 s 13434 2315 13542 2425 4 gnd
port 517 nsew
rlabel metal2 s 18426 21275 18534 21385 4 gnd
port 517 nsew
rlabel metal2 s 13434 9205 13542 9281 4 gnd
port 517 nsew
rlabel metal2 s 8922 9205 9030 9281 4 gnd
port 517 nsew
rlabel metal2 s 18906 20485 19014 20595 4 gnd
port 517 nsew
rlabel metal2 s 19674 20739 19782 20815 4 gnd
port 517 nsew
rlabel metal2 s 18906 12049 19014 12125 4 gnd
port 517 nsew
rlabel metal2 s 8922 7055 9030 7165 4 gnd
port 517 nsew
rlabel metal2 s 3450 3895 3558 4005 4 gnd
port 517 nsew
rlabel metal2 s 7194 15525 7302 15601 4 gnd
port 517 nsew
rlabel metal2 s 11418 22319 11526 22395 4 gnd
port 517 nsew
rlabel metal2 s 186 2095 294 2171 4 gnd
port 517 nsew
rlabel metal2 s 5946 5475 6054 5585 4 gnd
port 517 nsew
rlabel metal2 s 9690 5475 9798 5585 4 gnd
port 517 nsew
rlabel metal2 s 17178 11575 17286 11651 4 gnd
port 517 nsew
rlabel metal2 s 7194 15999 7302 16075 4 gnd
port 517 nsew
rlabel metal2 s 4698 9205 4806 9281 4 gnd
port 517 nsew
rlabel metal2 s 186 735 294 845 4 gnd
port 517 nsew
rlabel metal2 s 10170 22635 10278 22711 4 gnd
port 517 nsew
rlabel metal2 s 16410 19949 16518 20025 4 gnd
port 517 nsew
rlabel metal2 s 9690 17105 9798 17181 4 gnd
port 517 nsew
rlabel metal2 s 3930 9995 4038 10071 4 gnd
port 517 nsew
rlabel metal2 s 12186 14735 12294 14811 4 gnd
port 517 nsew
rlabel metal2 s 19674 -55 19782 55 4 gnd
port 517 nsew
rlabel metal2 s 6426 15745 6534 15855 4 gnd
port 517 nsew
rlabel metal2 s 7674 12839 7782 12915 4 gnd
port 517 nsew
rlabel metal2 s 12666 14735 12774 14811 4 gnd
port 517 nsew
rlabel metal2 s 954 3105 1062 3215 4 gnd
port 517 nsew
rlabel metal2 s 10170 3105 10278 3215 4 gnd
port 517 nsew
rlabel metal2 s 3930 16535 4038 16645 4 gnd
port 517 nsew
rlabel metal2 s 15162 4939 15270 5015 4 gnd
port 517 nsew
rlabel metal2 s 10938 17325 11046 17435 4 gnd
port 517 nsew
rlabel metal2 s 11418 18369 11526 18445 4 gnd
port 517 nsew
rlabel metal2 s 13914 3675 14022 3751 4 gnd
port 517 nsew
rlabel metal2 s 954 6045 1062 6121 4 gnd
port 517 nsew
rlabel metal2 s 7194 735 7302 845 4 gnd
port 517 nsew
rlabel metal2 s 17178 25005 17286 25081 4 gnd
port 517 nsew
rlabel metal2 s 5946 9205 6054 9281 4 gnd
port 517 nsew
rlabel metal2 s 3450 12839 3558 12915 4 gnd
port 517 nsew
rlabel metal2 s 11418 4939 11526 5015 4 gnd
port 517 nsew
rlabel metal2 s 10938 6519 11046 6595 4 gnd
port 517 nsew
rlabel metal2 s 10170 4939 10278 5015 4 gnd
port 517 nsew
rlabel metal2 s 954 19695 1062 19805 4 gnd
port 517 nsew
rlabel metal2 s 18426 11795 18534 11905 4 gnd
port 517 nsew
rlabel metal2 s 17178 25225 17286 25335 4 gnd
port 517 nsew
rlabel metal2 s 2202 19695 2310 19805 4 gnd
port 517 nsew
rlabel metal2 s 5178 8635 5286 8745 4 gnd
port 517 nsew
rlabel metal2 s 8442 14735 8550 14811 4 gnd
port 517 nsew
rlabel metal2 s 1434 5729 1542 5805 4 gnd
port 517 nsew
rlabel metal2 s 2682 12585 2790 12695 4 gnd
port 517 nsew
rlabel metal2 s 13434 10215 13542 10325 4 gnd
port 517 nsew
rlabel metal2 s 11418 5255 11526 5331 4 gnd
port 517 nsew
rlabel metal2 s 17178 10215 17286 10325 4 gnd
port 517 nsew
rlabel metal2 s 14682 3675 14790 3751 4 gnd
port 517 nsew
rlabel metal2 s 12186 16315 12294 16391 4 gnd
port 517 nsew
rlabel metal2 s 15930 21055 16038 21131 4 gnd
port 517 nsew
rlabel metal2 s 2202 15745 2310 15855 4 gnd
port 517 nsew
rlabel metal2 s 12186 17105 12294 17181 4 gnd
port 517 nsew
rlabel metal2 s 15930 10469 16038 10545 4 gnd
port 517 nsew
rlabel metal2 s 12186 23425 12294 23501 4 gnd
port 517 nsew
rlabel metal2 s 12666 16315 12774 16391 4 gnd
port 517 nsew
rlabel metal2 s 15930 22635 16038 22711 4 gnd
port 517 nsew
rlabel metal2 s 5946 16789 6054 16865 4 gnd
port 517 nsew
rlabel metal2 s 12666 4465 12774 4541 4 gnd
port 517 nsew
rlabel metal2 s 14682 12839 14790 12915 4 gnd
port 517 nsew
rlabel metal2 s 186 16315 294 16391 4 gnd
port 517 nsew
rlabel metal2 s 9690 15999 9798 16075 4 gnd
port 517 nsew
rlabel metal2 s 1434 14165 1542 14275 4 gnd
port 517 nsew
rlabel metal2 s 5178 8099 5286 8175 4 gnd
port 517 nsew
rlabel metal2 s 186 21845 294 21921 4 gnd
port 517 nsew
rlabel metal2 s 15930 10785 16038 10861 4 gnd
port 517 nsew
rlabel metal2 s 5178 11575 5286 11651 4 gnd
port 517 nsew
rlabel metal2 s 12186 23645 12294 23755 4 gnd
port 517 nsew
rlabel metal2 s 18426 4465 18534 4541 4 gnd
port 517 nsew
rlabel metal2 s 15162 19475 15270 19551 4 gnd
port 517 nsew
rlabel metal2 s 12186 7055 12294 7165 4 gnd
port 517 nsew
rlabel metal2 s 13434 9679 13542 9755 4 gnd
port 517 nsew
rlabel metal2 s 7194 3359 7302 3435 4 gnd
port 517 nsew
rlabel metal2 s 954 14735 1062 14811 4 gnd
port 517 nsew
rlabel metal2 s 4698 10215 4806 10325 4 gnd
port 517 nsew
rlabel metal2 s 12666 23109 12774 23185 4 gnd
port 517 nsew
rlabel metal2 s 18426 22635 18534 22711 4 gnd
port 517 nsew
rlabel metal2 s 9690 -55 9798 55 4 gnd
port 517 nsew
rlabel metal2 s 13434 5475 13542 5585 4 gnd
port 517 nsew
rlabel metal2 s 7674 3105 7782 3215 4 gnd
port 517 nsew
rlabel metal2 s 10170 19949 10278 20025 4 gnd
port 517 nsew
rlabel metal2 s 13914 13945 14022 14021 4 gnd
port 517 nsew
rlabel metal2 s 5178 2569 5286 2645 4 gnd
port 517 nsew
rlabel metal2 s 8442 989 8550 1065 4 gnd
port 517 nsew
rlabel metal2 s 2202 23109 2310 23185 4 gnd
port 517 nsew
rlabel metal2 s 14682 11259 14790 11335 4 gnd
port 517 nsew
rlabel metal2 s 5946 6835 6054 6911 4 gnd
port 517 nsew
rlabel metal2 s 186 5729 294 5805 4 gnd
port 517 nsew
rlabel metal2 s 2682 18115 2790 18225 4 gnd
port 517 nsew
rlabel metal2 s 13434 14165 13542 14275 4 gnd
port 517 nsew
rlabel metal2 s 18906 25005 19014 25081 4 gnd
port 517 nsew
rlabel metal2 s 18906 6835 19014 6911 4 gnd
port 517 nsew
rlabel metal2 s 2682 10215 2790 10325 4 gnd
port 517 nsew
rlabel metal2 s 7194 17105 7302 17181 4 gnd
port 517 nsew
rlabel metal2 s 7674 12049 7782 12125 4 gnd
port 517 nsew
rlabel metal2 s 954 14419 1062 14495 4 gnd
port 517 nsew
rlabel metal2 s 17178 14955 17286 15065 4 gnd
port 517 nsew
rlabel metal2 s 954 19159 1062 19235 4 gnd
port 517 nsew
rlabel metal2 s 12666 14165 12774 14275 4 gnd
port 517 nsew
rlabel metal2 s 17658 7845 17766 7955 4 gnd
port 517 nsew
rlabel metal2 s 4698 17325 4806 17435 4 gnd
port 517 nsew
rlabel metal2 s 10938 11259 11046 11335 4 gnd
port 517 nsew
rlabel metal2 s 12186 2885 12294 2961 4 gnd
port 517 nsew
rlabel metal2 s 9690 10215 9798 10325 4 gnd
port 517 nsew
rlabel metal2 s 17178 4685 17286 4795 4 gnd
port 517 nsew
rlabel metal2 s 9690 2315 9798 2425 4 gnd
port 517 nsew
rlabel metal2 s 12666 8635 12774 8745 4 gnd
port 517 nsew
rlabel metal2 s 13914 1305 14022 1381 4 gnd
port 517 nsew
rlabel metal2 s 16410 11795 16518 11905 4 gnd
port 517 nsew
rlabel metal2 s 10170 3359 10278 3435 4 gnd
port 517 nsew
rlabel metal2 s 10170 17105 10278 17181 4 gnd
port 517 nsew
rlabel metal2 s 12666 20739 12774 20815 4 gnd
port 517 nsew
rlabel metal2 s 3450 21055 3558 21131 4 gnd
port 517 nsew
rlabel metal2 s 1434 22319 1542 22395 4 gnd
port 517 nsew
rlabel metal2 s 954 23645 1062 23755 4 gnd
port 517 nsew
rlabel metal2 s 2682 18369 2790 18445 4 gnd
port 517 nsew
rlabel metal2 s 5178 24215 5286 24291 4 gnd
port 517 nsew
rlabel metal2 s 14682 19695 14790 19805 4 gnd
port 517 nsew
rlabel metal2 s 954 21845 1062 21921 4 gnd
port 517 nsew
rlabel metal2 s 7194 18369 7302 18445 4 gnd
port 517 nsew
rlabel metal2 s 15162 15999 15270 16075 4 gnd
port 517 nsew
rlabel metal2 s 10170 22319 10278 22395 4 gnd
port 517 nsew
rlabel metal2 s 2202 24435 2310 24545 4 gnd
port 517 nsew
rlabel metal2 s 19674 11795 19782 11905 4 gnd
port 517 nsew
rlabel metal2 s 5178 13155 5286 13231 4 gnd
port 517 nsew
rlabel metal2 s 2202 7055 2310 7165 4 gnd
port 517 nsew
rlabel metal2 s 3930 7055 4038 7165 4 gnd
port 517 nsew
rlabel metal2 s 13914 22635 14022 22711 4 gnd
port 517 nsew
rlabel metal2 s 6426 3105 6534 3215 4 gnd
port 517 nsew
rlabel metal2 s 9690 199 9798 275 4 gnd
port 517 nsew
rlabel metal2 s 10170 4685 10278 4795 4 gnd
port 517 nsew
rlabel metal2 s 18426 9995 18534 10071 4 gnd
port 517 nsew
rlabel metal2 s 14682 19159 14790 19235 4 gnd
port 517 nsew
rlabel metal2 s 15930 19475 16038 19551 4 gnd
port 517 nsew
rlabel metal2 s 7674 3895 7782 4005 4 gnd
port 517 nsew
rlabel metal2 s 186 22065 294 22175 4 gnd
port 517 nsew
rlabel metal2 s 2682 24215 2790 24291 4 gnd
port 517 nsew
rlabel metal2 s 15162 4685 15270 4795 4 gnd
port 517 nsew
rlabel metal2 s 12186 17325 12294 17435 4 gnd
port 517 nsew
rlabel metal2 s 12186 17895 12294 17971 4 gnd
port 517 nsew
rlabel metal2 s 9690 2885 9798 2961 4 gnd
port 517 nsew
rlabel metal2 s 8442 9425 8550 9535 4 gnd
port 517 nsew
rlabel metal2 s 8442 8889 8550 8965 4 gnd
port 517 nsew
rlabel metal2 s 1434 11575 1542 11651 4 gnd
port 517 nsew
rlabel metal2 s 954 12585 1062 12695 4 gnd
port 517 nsew
rlabel metal2 s 2202 8415 2310 8491 4 gnd
port 517 nsew
rlabel metal2 s 15162 21845 15270 21921 4 gnd
port 517 nsew
rlabel metal2 s 18426 14165 18534 14275 4 gnd
port 517 nsew
rlabel metal2 s 19674 2315 19782 2425 4 gnd
port 517 nsew
rlabel metal2 s 15162 8099 15270 8175 4 gnd
port 517 nsew
rlabel metal2 s 11418 13945 11526 14021 4 gnd
port 517 nsew
rlabel metal2 s 11418 10785 11526 10861 4 gnd
port 517 nsew
rlabel metal2 s 18426 2095 18534 2171 4 gnd
port 517 nsew
rlabel metal2 s 12666 2095 12774 2171 4 gnd
port 517 nsew
rlabel metal2 s 7674 2569 7782 2645 4 gnd
port 517 nsew
rlabel metal2 s 7194 21529 7302 21605 4 gnd
port 517 nsew
rlabel metal2 s 4698 12585 4806 12695 4 gnd
port 517 nsew
rlabel metal2 s 12186 6835 12294 6911 4 gnd
port 517 nsew
rlabel metal2 s 9690 24689 9798 24765 4 gnd
port 517 nsew
rlabel metal2 s 10938 11005 11046 11115 4 gnd
port 517 nsew
rlabel metal2 s 5178 16789 5286 16865 4 gnd
port 517 nsew
rlabel metal2 s 14682 15525 14790 15601 4 gnd
port 517 nsew
rlabel metal2 s 5946 22319 6054 22395 4 gnd
port 517 nsew
rlabel metal2 s 7194 24435 7302 24545 4 gnd
port 517 nsew
rlabel metal2 s 15930 21845 16038 21921 4 gnd
port 517 nsew
rlabel metal2 s 5946 24215 6054 24291 4 gnd
port 517 nsew
rlabel metal2 s 186 8099 294 8175 4 gnd
port 517 nsew
rlabel metal2 s 19674 7625 19782 7701 4 gnd
port 517 nsew
rlabel metal2 s 12666 7309 12774 7385 4 gnd
port 517 nsew
rlabel metal2 s 18426 3895 18534 4005 4 gnd
port 517 nsew
rlabel metal2 s 19674 22635 19782 22711 4 gnd
port 517 nsew
rlabel metal2 s 2682 3895 2790 4005 4 gnd
port 517 nsew
rlabel metal2 s 5178 14735 5286 14811 4 gnd
port 517 nsew
rlabel metal2 s 10170 22855 10278 22965 4 gnd
port 517 nsew
rlabel metal2 s 12666 12585 12774 12695 4 gnd
port 517 nsew
rlabel metal2 s 15162 8889 15270 8965 4 gnd
port 517 nsew
rlabel metal2 s 18906 11259 19014 11335 4 gnd
port 517 nsew
rlabel metal2 s 17178 18685 17286 18761 4 gnd
port 517 nsew
rlabel metal2 s 4698 22319 4806 22395 4 gnd
port 517 nsew
rlabel metal2 s 3930 18115 4038 18225 4 gnd
port 517 nsew
rlabel metal2 s 13434 3895 13542 4005 4 gnd
port 517 nsew
rlabel metal2 s 15930 3105 16038 3215 4 gnd
port 517 nsew
rlabel metal2 s 14682 13945 14790 14021 4 gnd
port 517 nsew
rlabel metal2 s 4698 12049 4806 12125 4 gnd
port 517 nsew
rlabel metal2 s 186 7309 294 7385 4 gnd
port 517 nsew
rlabel metal2 s 5946 6519 6054 6595 4 gnd
port 517 nsew
rlabel metal2 s 9690 5255 9798 5331 4 gnd
port 517 nsew
rlabel metal2 s 3930 20265 4038 20341 4 gnd
port 517 nsew
rlabel metal2 s 4698 18115 4806 18225 4 gnd
port 517 nsew
rlabel metal2 s 1434 24689 1542 24765 4 gnd
port 517 nsew
rlabel metal2 s 9690 15209 9798 15285 4 gnd
port 517 nsew
rlabel metal2 s 954 13629 1062 13705 4 gnd
port 517 nsew
rlabel metal2 s 14682 22319 14790 22395 4 gnd
port 517 nsew
rlabel metal2 s 15162 20485 15270 20595 4 gnd
port 517 nsew
rlabel metal2 s 2682 6519 2790 6595 4 gnd
port 517 nsew
rlabel metal2 s 15930 2315 16038 2425 4 gnd
port 517 nsew
rlabel metal2 s 12666 24435 12774 24545 4 gnd
port 517 nsew
rlabel metal2 s 13914 7845 14022 7955 4 gnd
port 517 nsew
rlabel metal2 s 13914 21529 14022 21605 4 gnd
port 517 nsew
rlabel metal2 s 8442 9205 8550 9281 4 gnd
port 517 nsew
rlabel metal2 s 2682 18685 2790 18761 4 gnd
port 517 nsew
rlabel metal2 s 954 23109 1062 23185 4 gnd
port 517 nsew
rlabel metal2 s 12186 10469 12294 10545 4 gnd
port 517 nsew
rlabel metal2 s 7194 12839 7302 12915 4 gnd
port 517 nsew
rlabel metal2 s 9690 989 9798 1065 4 gnd
port 517 nsew
rlabel metal2 s 11418 15999 11526 16075 4 gnd
port 517 nsew
rlabel metal2 s 7194 12365 7302 12441 4 gnd
port 517 nsew
rlabel metal2 s 13434 13945 13542 14021 4 gnd
port 517 nsew
rlabel metal2 s 5178 18905 5286 19015 4 gnd
port 517 nsew
rlabel metal2 s 19674 8889 19782 8965 4 gnd
port 517 nsew
rlabel metal2 s 7674 14419 7782 14495 4 gnd
port 517 nsew
rlabel metal2 s 2202 25005 2310 25081 4 gnd
port 517 nsew
rlabel metal2 s 186 -55 294 55 4 gnd
port 517 nsew
rlabel metal2 s 7674 9205 7782 9281 4 gnd
port 517 nsew
rlabel metal2 s 12186 9425 12294 9535 4 gnd
port 517 nsew
rlabel metal2 s 3450 17325 3558 17435 4 gnd
port 517 nsew
rlabel metal2 s 8442 11795 8550 11905 4 gnd
port 517 nsew
rlabel metal2 s 954 6835 1062 6911 4 gnd
port 517 nsew
rlabel metal2 s 8922 7309 9030 7385 4 gnd
port 517 nsew
rlabel metal2 s 13434 17105 13542 17181 4 gnd
port 517 nsew
rlabel metal2 s 15162 17325 15270 17435 4 gnd
port 517 nsew
rlabel metal2 s 3930 5729 4038 5805 4 gnd
port 517 nsew
rlabel metal2 s 2682 22319 2790 22395 4 gnd
port 517 nsew
rlabel metal2 s 13434 13155 13542 13231 4 gnd
port 517 nsew
rlabel metal2 s 10938 14735 11046 14811 4 gnd
port 517 nsew
rlabel metal2 s 2202 3895 2310 4005 4 gnd
port 517 nsew
rlabel metal2 s 11418 3105 11526 3215 4 gnd
port 517 nsew
rlabel metal2 s 5946 19475 6054 19551 4 gnd
port 517 nsew
rlabel metal2 s 8922 21055 9030 21131 4 gnd
port 517 nsew
rlabel metal2 s 3930 13629 4038 13705 4 gnd
port 517 nsew
rlabel metal2 s 11418 8099 11526 8175 4 gnd
port 517 nsew
rlabel metal2 s 1434 11005 1542 11115 4 gnd
port 517 nsew
rlabel metal2 s 2682 20485 2790 20595 4 gnd
port 517 nsew
rlabel metal2 s 7674 11005 7782 11115 4 gnd
port 517 nsew
rlabel metal2 s 5946 2095 6054 2171 4 gnd
port 517 nsew
rlabel metal2 s 15930 24689 16038 24765 4 gnd
port 517 nsew
rlabel metal2 s 16410 10469 16518 10545 4 gnd
port 517 nsew
rlabel metal2 s 10170 11575 10278 11651 4 gnd
port 517 nsew
rlabel metal2 s 12186 12365 12294 12441 4 gnd
port 517 nsew
rlabel metal2 s 12666 20485 12774 20595 4 gnd
port 517 nsew
rlabel metal2 s 13914 13375 14022 13485 4 gnd
port 517 nsew
rlabel metal2 s 954 21275 1062 21385 4 gnd
port 517 nsew
rlabel metal2 s 4698 9425 4806 9535 4 gnd
port 517 nsew
rlabel metal2 s 11418 21275 11526 21385 4 gnd
port 517 nsew
rlabel metal2 s 10170 16789 10278 16865 4 gnd
port 517 nsew
rlabel metal2 s 17178 17579 17286 17655 4 gnd
port 517 nsew
rlabel metal2 s 13914 11259 14022 11335 4 gnd
port 517 nsew
rlabel metal2 s 186 25225 294 25335 4 gnd
port 517 nsew
rlabel metal2 s 18426 8635 18534 8745 4 gnd
port 517 nsew
rlabel metal2 s 3930 735 4038 845 4 gnd
port 517 nsew
rlabel metal2 s 18906 1305 19014 1381 4 gnd
port 517 nsew
rlabel metal2 s 17658 14419 17766 14495 4 gnd
port 517 nsew
rlabel metal2 s 17658 1779 17766 1855 4 gnd
port 517 nsew
rlabel metal2 s 6426 23109 6534 23185 4 gnd
port 517 nsew
rlabel metal2 s 5178 735 5286 845 4 gnd
port 517 nsew
rlabel metal2 s 7674 8635 7782 8745 4 gnd
port 517 nsew
rlabel metal2 s 14682 13155 14790 13231 4 gnd
port 517 nsew
rlabel metal2 s 19674 22855 19782 22965 4 gnd
port 517 nsew
rlabel metal2 s 7674 1305 7782 1381 4 gnd
port 517 nsew
rlabel metal2 s 16410 6519 16518 6595 4 gnd
port 517 nsew
rlabel metal2 s 2202 16535 2310 16645 4 gnd
port 517 nsew
rlabel metal2 s 8442 16315 8550 16391 4 gnd
port 517 nsew
rlabel metal2 s 13914 24215 14022 24291 4 gnd
port 517 nsew
rlabel metal2 s 3450 8635 3558 8745 4 gnd
port 517 nsew
rlabel metal2 s 2682 7845 2790 7955 4 gnd
port 517 nsew
rlabel metal2 s 186 7845 294 7955 4 gnd
port 517 nsew
rlabel metal2 s 9690 14419 9798 14495 4 gnd
port 517 nsew
rlabel metal2 s 7194 22855 7302 22965 4 gnd
port 517 nsew
rlabel metal2 s 954 6519 1062 6595 4 gnd
port 517 nsew
rlabel metal2 s 13914 1779 14022 1855 4 gnd
port 517 nsew
rlabel metal2 s 11418 7625 11526 7701 4 gnd
port 517 nsew
rlabel metal2 s 11418 21529 11526 21605 4 gnd
port 517 nsew
rlabel metal2 s 19674 2569 19782 2645 4 gnd
port 517 nsew
rlabel metal2 s 186 8889 294 8965 4 gnd
port 517 nsew
rlabel metal2 s 13914 9425 14022 9535 4 gnd
port 517 nsew
rlabel metal2 s 14682 10469 14790 10545 4 gnd
port 517 nsew
rlabel metal2 s 2202 4685 2310 4795 4 gnd
port 517 nsew
rlabel metal2 s 2202 12839 2310 12915 4 gnd
port 517 nsew
rlabel metal2 s 5946 9425 6054 9535 4 gnd
port 517 nsew
rlabel metal2 s 1434 20485 1542 20595 4 gnd
port 517 nsew
rlabel metal2 s 11418 15525 11526 15601 4 gnd
port 517 nsew
rlabel metal2 s 4698 6519 4806 6595 4 gnd
port 517 nsew
rlabel metal2 s 2202 -55 2310 55 4 gnd
port 517 nsew
rlabel metal2 s 8442 3359 8550 3435 4 gnd
port 517 nsew
rlabel metal2 s 8442 18369 8550 18445 4 gnd
port 517 nsew
rlabel metal2 s 17658 13629 17766 13705 4 gnd
port 517 nsew
rlabel metal2 s 18906 17895 19014 17971 4 gnd
port 517 nsew
rlabel metal2 s 5946 22635 6054 22711 4 gnd
port 517 nsew
rlabel metal2 s 186 13155 294 13231 4 gnd
port 517 nsew
rlabel metal2 s 10170 14735 10278 14811 4 gnd
port 517 nsew
rlabel metal2 s 10170 6519 10278 6595 4 gnd
port 517 nsew
rlabel metal2 s 12666 4149 12774 4225 4 gnd
port 517 nsew
rlabel metal2 s 3450 21529 3558 21605 4 gnd
port 517 nsew
rlabel metal2 s 15930 17579 16038 17655 4 gnd
port 517 nsew
rlabel metal2 s 6426 4939 6534 5015 4 gnd
port 517 nsew
rlabel metal2 s 18426 13375 18534 13485 4 gnd
port 517 nsew
rlabel metal2 s 8922 15209 9030 15285 4 gnd
port 517 nsew
rlabel metal2 s 5946 6045 6054 6121 4 gnd
port 517 nsew
rlabel metal2 s 954 3359 1062 3435 4 gnd
port 517 nsew
rlabel metal2 s 14682 24215 14790 24291 4 gnd
port 517 nsew
rlabel metal2 s 15162 735 15270 845 4 gnd
port 517 nsew
rlabel metal2 s 6426 4149 6534 4225 4 gnd
port 517 nsew
rlabel metal2 s 18906 23899 19014 23975 4 gnd
port 517 nsew
rlabel metal2 s 12186 8635 12294 8745 4 gnd
port 517 nsew
rlabel metal2 s 12186 23109 12294 23185 4 gnd
port 517 nsew
rlabel metal2 s 10938 25005 11046 25081 4 gnd
port 517 nsew
rlabel metal2 s 3450 25005 3558 25081 4 gnd
port 517 nsew
rlabel metal2 s 8922 515 9030 591 4 gnd
port 517 nsew
rlabel metal2 s 17178 8099 17286 8175 4 gnd
port 517 nsew
rlabel metal2 s 954 22635 1062 22711 4 gnd
port 517 nsew
rlabel metal2 s 12666 22635 12774 22711 4 gnd
port 517 nsew
rlabel metal2 s 12186 515 12294 591 4 gnd
port 517 nsew
rlabel metal2 s 15930 6519 16038 6595 4 gnd
port 517 nsew
rlabel metal2 s 8922 25225 9030 25335 4 gnd
port 517 nsew
rlabel metal2 s 2682 20265 2790 20341 4 gnd
port 517 nsew
rlabel metal2 s 7194 18905 7302 19015 4 gnd
port 517 nsew
rlabel metal2 s 16410 19159 16518 19235 4 gnd
port 517 nsew
rlabel metal2 s 13434 7055 13542 7165 4 gnd
port 517 nsew
rlabel metal2 s 10938 7625 11046 7701 4 gnd
port 517 nsew
rlabel metal2 s 13434 12365 13542 12441 4 gnd
port 517 nsew
rlabel metal2 s 18426 17579 18534 17655 4 gnd
port 517 nsew
rlabel metal2 s 2682 11005 2790 11115 4 gnd
port 517 nsew
rlabel metal2 s 10938 7055 11046 7165 4 gnd
port 517 nsew
rlabel metal2 s 17178 17105 17286 17181 4 gnd
port 517 nsew
rlabel metal2 s 954 22855 1062 22965 4 gnd
port 517 nsew
rlabel metal2 s 2682 11575 2790 11651 4 gnd
port 517 nsew
rlabel metal2 s 3930 4939 4038 5015 4 gnd
port 517 nsew
rlabel metal2 s 7194 22319 7302 22395 4 gnd
port 517 nsew
rlabel metal2 s 9690 1525 9798 1635 4 gnd
port 517 nsew
rlabel metal2 s 16410 8099 16518 8175 4 gnd
port 517 nsew
rlabel metal2 s 10170 12365 10278 12441 4 gnd
port 517 nsew
rlabel metal2 s 1434 20739 1542 20815 4 gnd
port 517 nsew
rlabel metal2 s 14682 4149 14790 4225 4 gnd
port 517 nsew
rlabel metal2 s 7194 17895 7302 17971 4 gnd
port 517 nsew
rlabel metal2 s 15930 23425 16038 23501 4 gnd
port 517 nsew
rlabel metal2 s 15930 16535 16038 16645 4 gnd
port 517 nsew
rlabel metal2 s 13434 19949 13542 20025 4 gnd
port 517 nsew
rlabel metal2 s 15930 199 16038 275 4 gnd
port 517 nsew
rlabel metal2 s 5178 15745 5286 15855 4 gnd
port 517 nsew
rlabel metal2 s 10938 9995 11046 10071 4 gnd
port 517 nsew
rlabel metal2 s 15930 15209 16038 15285 4 gnd
port 517 nsew
rlabel metal2 s 4698 13155 4806 13231 4 gnd
port 517 nsew
rlabel metal2 s 7674 6265 7782 6375 4 gnd
port 517 nsew
rlabel metal2 s 1434 7625 1542 7701 4 gnd
port 517 nsew
rlabel metal2 s 5946 8099 6054 8175 4 gnd
port 517 nsew
rlabel metal2 s 5178 13375 5286 13485 4 gnd
port 517 nsew
rlabel metal2 s 13914 11005 14022 11115 4 gnd
port 517 nsew
rlabel metal2 s 17178 20485 17286 20595 4 gnd
port 517 nsew
rlabel metal2 s 11418 -55 11526 55 4 gnd
port 517 nsew
rlabel metal2 s 4698 17895 4806 17971 4 gnd
port 517 nsew
rlabel metal2 s 6426 2569 6534 2645 4 gnd
port 517 nsew
rlabel metal2 s 18906 515 19014 591 4 gnd
port 517 nsew
rlabel metal2 s 17658 2885 17766 2961 4 gnd
port 517 nsew
rlabel metal2 s 954 5255 1062 5331 4 gnd
port 517 nsew
rlabel metal2 s 10170 11795 10278 11905 4 gnd
port 517 nsew
rlabel metal2 s 7194 18115 7302 18225 4 gnd
port 517 nsew
rlabel metal2 s 17178 8415 17286 8491 4 gnd
port 517 nsew
rlabel metal2 s 17658 10215 17766 10325 4 gnd
port 517 nsew
rlabel metal2 s 18906 20739 19014 20815 4 gnd
port 517 nsew
rlabel metal2 s 19674 10785 19782 10861 4 gnd
port 517 nsew
rlabel metal2 s 6426 3359 6534 3435 4 gnd
port 517 nsew
rlabel metal2 s 12666 8415 12774 8491 4 gnd
port 517 nsew
rlabel metal2 s 18906 18685 19014 18761 4 gnd
port 517 nsew
rlabel metal2 s 19674 23645 19782 23755 4 gnd
port 517 nsew
rlabel metal2 s 19674 9679 19782 9755 4 gnd
port 517 nsew
rlabel metal2 s 16410 9679 16518 9755 4 gnd
port 517 nsew
rlabel metal2 s 8442 2095 8550 2171 4 gnd
port 517 nsew
rlabel metal2 s 6426 5255 6534 5331 4 gnd
port 517 nsew
rlabel metal2 s 8442 23425 8550 23501 4 gnd
port 517 nsew
rlabel metal2 s 18426 24215 18534 24291 4 gnd
port 517 nsew
rlabel metal2 s 13914 12839 14022 12915 4 gnd
port 517 nsew
rlabel metal2 s 9690 7625 9798 7701 4 gnd
port 517 nsew
rlabel metal2 s 5178 4685 5286 4795 4 gnd
port 517 nsew
rlabel metal2 s 13434 20265 13542 20341 4 gnd
port 517 nsew
rlabel metal2 s 10170 6265 10278 6375 4 gnd
port 517 nsew
rlabel metal2 s 11418 24435 11526 24545 4 gnd
port 517 nsew
rlabel metal2 s 17658 19695 17766 19805 4 gnd
port 517 nsew
rlabel metal2 s 13434 19159 13542 19235 4 gnd
port 517 nsew
rlabel metal2 s 4698 18905 4806 19015 4 gnd
port 517 nsew
rlabel metal2 s 2202 13375 2310 13485 4 gnd
port 517 nsew
rlabel metal2 s 6426 22635 6534 22711 4 gnd
port 517 nsew
rlabel metal2 s 11418 14955 11526 15065 4 gnd
port 517 nsew
rlabel metal2 s 3930 17895 4038 17971 4 gnd
port 517 nsew
rlabel metal2 s 17178 8635 17286 8745 4 gnd
port 517 nsew
rlabel metal2 s 17658 13945 17766 14021 4 gnd
port 517 nsew
rlabel metal2 s 10938 2569 11046 2645 4 gnd
port 517 nsew
rlabel metal2 s 5946 -55 6054 55 4 gnd
port 517 nsew
rlabel metal2 s 2682 9425 2790 9535 4 gnd
port 517 nsew
rlabel metal2 s 6426 18115 6534 18225 4 gnd
port 517 nsew
rlabel metal2 s 16410 25005 16518 25081 4 gnd
port 517 nsew
rlabel metal2 s 17178 5729 17286 5805 4 gnd
port 517 nsew
rlabel metal2 s 1434 19159 1542 19235 4 gnd
port 517 nsew
rlabel metal2 s 954 13945 1062 14021 4 gnd
port 517 nsew
rlabel metal2 s 2202 24215 2310 24291 4 gnd
port 517 nsew
rlabel metal2 s 6426 20485 6534 20595 4 gnd
port 517 nsew
rlabel metal2 s 10938 4465 11046 4541 4 gnd
port 517 nsew
rlabel metal2 s 15162 18685 15270 18761 4 gnd
port 517 nsew
rlabel metal2 s 5946 12839 6054 12915 4 gnd
port 517 nsew
rlabel metal2 s 2202 14955 2310 15065 4 gnd
port 517 nsew
rlabel metal2 s 3930 8415 4038 8491 4 gnd
port 517 nsew
rlabel metal2 s 3930 21529 4038 21605 4 gnd
port 517 nsew
rlabel metal2 s 11418 11005 11526 11115 4 gnd
port 517 nsew
rlabel metal2 s 186 5475 294 5585 4 gnd
port 517 nsew
rlabel metal2 s 10938 19159 11046 19235 4 gnd
port 517 nsew
rlabel metal2 s 3930 2569 4038 2645 4 gnd
port 517 nsew
rlabel metal2 s 11418 1779 11526 1855 4 gnd
port 517 nsew
rlabel metal2 s 12186 14419 12294 14495 4 gnd
port 517 nsew
rlabel metal2 s 13434 11795 13542 11905 4 gnd
port 517 nsew
rlabel metal2 s 13434 12839 13542 12915 4 gnd
port 517 nsew
rlabel metal2 s 18906 16315 19014 16391 4 gnd
port 517 nsew
rlabel metal2 s 17178 6265 17286 6375 4 gnd
port 517 nsew
rlabel metal2 s 11418 7055 11526 7165 4 gnd
port 517 nsew
rlabel metal2 s 7194 10469 7302 10545 4 gnd
port 517 nsew
rlabel metal2 s 16410 22855 16518 22965 4 gnd
port 517 nsew
rlabel metal2 s 15930 7309 16038 7385 4 gnd
port 517 nsew
rlabel metal2 s 18906 23645 19014 23755 4 gnd
port 517 nsew
rlabel metal2 s 19674 8415 19782 8491 4 gnd
port 517 nsew
rlabel metal2 s 7194 13155 7302 13231 4 gnd
port 517 nsew
rlabel metal2 s 2682 15209 2790 15285 4 gnd
port 517 nsew
rlabel metal2 s 17658 9995 17766 10071 4 gnd
port 517 nsew
rlabel metal2 s 5946 18115 6054 18225 4 gnd
port 517 nsew
rlabel metal2 s 18906 9679 19014 9755 4 gnd
port 517 nsew
rlabel metal2 s 10170 18905 10278 19015 4 gnd
port 517 nsew
rlabel metal2 s 9690 9995 9798 10071 4 gnd
port 517 nsew
rlabel metal2 s 14682 1779 14790 1855 4 gnd
port 517 nsew
rlabel metal2 s 14682 17895 14790 17971 4 gnd
port 517 nsew
rlabel metal2 s 15930 15745 16038 15855 4 gnd
port 517 nsew
rlabel metal2 s 9690 1779 9798 1855 4 gnd
port 517 nsew
rlabel metal2 s 19674 1525 19782 1635 4 gnd
port 517 nsew
rlabel metal2 s 10170 24689 10278 24765 4 gnd
port 517 nsew
rlabel metal2 s 2202 4465 2310 4541 4 gnd
port 517 nsew
rlabel metal2 s 3450 9425 3558 9535 4 gnd
port 517 nsew
rlabel metal2 s 10938 15209 11046 15285 4 gnd
port 517 nsew
rlabel metal2 s 16410 6045 16518 6121 4 gnd
port 517 nsew
rlabel metal2 s 3930 23645 4038 23755 4 gnd
port 517 nsew
rlabel metal2 s 17178 735 17286 845 4 gnd
port 517 nsew
rlabel metal2 s 954 15525 1062 15601 4 gnd
port 517 nsew
rlabel metal2 s 7674 23425 7782 23501 4 gnd
port 517 nsew
rlabel metal2 s 13914 23425 14022 23501 4 gnd
port 517 nsew
rlabel metal2 s 2682 21055 2790 21131 4 gnd
port 517 nsew
rlabel metal2 s 10170 20265 10278 20341 4 gnd
port 517 nsew
rlabel metal2 s 19674 989 19782 1065 4 gnd
port 517 nsew
rlabel metal2 s 13914 11795 14022 11905 4 gnd
port 517 nsew
rlabel metal2 s 12186 22319 12294 22395 4 gnd
port 517 nsew
rlabel metal2 s 7674 11259 7782 11335 4 gnd
port 517 nsew
rlabel metal2 s 6426 18685 6534 18761 4 gnd
port 517 nsew
rlabel metal2 s 10938 20485 11046 20595 4 gnd
port 517 nsew
rlabel metal2 s 18906 18905 19014 19015 4 gnd
port 517 nsew
rlabel metal2 s 8922 2315 9030 2425 4 gnd
port 517 nsew
rlabel metal2 s 16410 3359 16518 3435 4 gnd
port 517 nsew
rlabel metal2 s 2202 6265 2310 6375 4 gnd
port 517 nsew
rlabel metal2 s 13434 22855 13542 22965 4 gnd
port 517 nsew
rlabel metal2 s 16410 11259 16518 11335 4 gnd
port 517 nsew
rlabel metal2 s 2202 25225 2310 25335 4 gnd
port 517 nsew
rlabel metal2 s 16410 23899 16518 23975 4 gnd
port 517 nsew
rlabel metal2 s 18426 23645 18534 23755 4 gnd
port 517 nsew
rlabel metal2 s 10170 3895 10278 4005 4 gnd
port 517 nsew
rlabel metal2 s 954 18685 1062 18761 4 gnd
port 517 nsew
rlabel metal2 s 2682 12839 2790 12915 4 gnd
port 517 nsew
rlabel metal2 s 13914 19475 14022 19551 4 gnd
port 517 nsew
rlabel metal2 s 13434 6835 13542 6911 4 gnd
port 517 nsew
rlabel metal2 s 2202 12365 2310 12441 4 gnd
port 517 nsew
rlabel metal2 s 2682 3675 2790 3751 4 gnd
port 517 nsew
rlabel metal2 s 18426 5475 18534 5585 4 gnd
port 517 nsew
rlabel metal2 s 3930 24435 4038 24545 4 gnd
port 517 nsew
rlabel metal2 s 5178 13629 5286 13705 4 gnd
port 517 nsew
rlabel metal2 s 13914 2095 14022 2171 4 gnd
port 517 nsew
rlabel metal2 s 17658 6835 17766 6911 4 gnd
port 517 nsew
rlabel metal2 s 17658 17579 17766 17655 4 gnd
port 517 nsew
rlabel metal2 s 3450 24215 3558 24291 4 gnd
port 517 nsew
rlabel metal2 s 9690 16315 9798 16391 4 gnd
port 517 nsew
rlabel metal2 s 12666 17105 12774 17181 4 gnd
port 517 nsew
rlabel metal2 s 19674 22319 19782 22395 4 gnd
port 517 nsew
rlabel metal2 s 9690 14955 9798 15065 4 gnd
port 517 nsew
rlabel metal2 s 5946 24689 6054 24765 4 gnd
port 517 nsew
rlabel metal2 s 1434 14735 1542 14811 4 gnd
port 517 nsew
rlabel metal2 s 7194 21275 7302 21385 4 gnd
port 517 nsew
rlabel metal2 s 8922 13629 9030 13705 4 gnd
port 517 nsew
rlabel metal2 s 19674 23425 19782 23501 4 gnd
port 517 nsew
rlabel metal2 s 8922 8635 9030 8745 4 gnd
port 517 nsew
rlabel metal2 s 7194 6519 7302 6595 4 gnd
port 517 nsew
rlabel metal2 s 3930 14735 4038 14811 4 gnd
port 517 nsew
rlabel metal2 s 2682 25005 2790 25081 4 gnd
port 517 nsew
rlabel metal2 s 8922 24435 9030 24545 4 gnd
port 517 nsew
rlabel metal2 s 7674 23109 7782 23185 4 gnd
port 517 nsew
rlabel metal2 s 4698 19159 4806 19235 4 gnd
port 517 nsew
rlabel metal2 s 9690 7845 9798 7955 4 gnd
port 517 nsew
rlabel metal2 s 5178 9679 5286 9755 4 gnd
port 517 nsew
rlabel metal2 s 15162 -55 15270 55 4 gnd
port 517 nsew
rlabel metal2 s 6426 17895 6534 17971 4 gnd
port 517 nsew
rlabel metal2 s 15930 1525 16038 1635 4 gnd
port 517 nsew
rlabel metal2 s 19674 24435 19782 24545 4 gnd
port 517 nsew
rlabel metal2 s 7674 21055 7782 21131 4 gnd
port 517 nsew
rlabel metal2 s 8442 199 8550 275 4 gnd
port 517 nsew
rlabel metal2 s 3450 17579 3558 17655 4 gnd
port 517 nsew
rlabel metal2 s 15930 18905 16038 19015 4 gnd
port 517 nsew
rlabel metal2 s 5946 21529 6054 21605 4 gnd
port 517 nsew
rlabel metal2 s 4698 7055 4806 7165 4 gnd
port 517 nsew
rlabel metal2 s 14682 13629 14790 13705 4 gnd
port 517 nsew
rlabel metal2 s 11418 7845 11526 7955 4 gnd
port 517 nsew
rlabel metal2 s 11418 12839 11526 12915 4 gnd
port 517 nsew
rlabel metal2 s 18906 7625 19014 7701 4 gnd
port 517 nsew
rlabel metal2 s 8922 -55 9030 55 4 gnd
port 517 nsew
rlabel metal2 s 13434 12585 13542 12695 4 gnd
port 517 nsew
rlabel metal2 s 18906 15999 19014 16075 4 gnd
port 517 nsew
rlabel metal2 s 19674 18905 19782 19015 4 gnd
port 517 nsew
rlabel metal2 s 2682 2315 2790 2425 4 gnd
port 517 nsew
rlabel metal2 s 16410 2095 16518 2171 4 gnd
port 517 nsew
rlabel metal2 s 17178 13375 17286 13485 4 gnd
port 517 nsew
rlabel metal2 s 18426 25005 18534 25081 4 gnd
port 517 nsew
rlabel metal2 s 2202 16789 2310 16865 4 gnd
port 517 nsew
rlabel metal2 s 14682 2095 14790 2171 4 gnd
port 517 nsew
rlabel metal2 s 19674 4939 19782 5015 4 gnd
port 517 nsew
rlabel metal2 s 16410 1525 16518 1635 4 gnd
port 517 nsew
rlabel metal2 s 3930 3675 4038 3751 4 gnd
port 517 nsew
rlabel metal2 s 7674 199 7782 275 4 gnd
port 517 nsew
rlabel metal2 s 18906 4685 19014 4795 4 gnd
port 517 nsew
rlabel metal2 s 14682 19475 14790 19551 4 gnd
port 517 nsew
rlabel metal2 s 8922 18905 9030 19015 4 gnd
port 517 nsew
rlabel metal2 s 13434 23109 13542 23185 4 gnd
port 517 nsew
rlabel metal2 s 5946 1305 6054 1381 4 gnd
port 517 nsew
rlabel metal2 s 12186 20485 12294 20595 4 gnd
port 517 nsew
rlabel metal2 s 3450 20265 3558 20341 4 gnd
port 517 nsew
rlabel metal2 s 12666 8889 12774 8965 4 gnd
port 517 nsew
rlabel metal2 s 8922 11005 9030 11115 4 gnd
port 517 nsew
rlabel metal2 s 2682 1779 2790 1855 4 gnd
port 517 nsew
rlabel metal2 s 17658 1525 17766 1635 4 gnd
port 517 nsew
rlabel metal2 s 17658 7309 17766 7385 4 gnd
port 517 nsew
rlabel metal2 s 3450 10785 3558 10861 4 gnd
port 517 nsew
rlabel metal2 s 6426 9679 6534 9755 4 gnd
port 517 nsew
rlabel metal2 s 17658 2315 17766 2425 4 gnd
port 517 nsew
rlabel metal2 s 18426 16789 18534 16865 4 gnd
port 517 nsew
rlabel metal2 s 15162 25225 15270 25335 4 gnd
port 517 nsew
rlabel metal2 s 13434 9995 13542 10071 4 gnd
port 517 nsew
rlabel metal2 s 8442 4465 8550 4541 4 gnd
port 517 nsew
rlabel metal2 s 4698 8415 4806 8491 4 gnd
port 517 nsew
rlabel metal2 s 18906 19695 19014 19805 4 gnd
port 517 nsew
rlabel metal2 s 12186 6045 12294 6121 4 gnd
port 517 nsew
rlabel metal2 s 18426 23899 18534 23975 4 gnd
port 517 nsew
rlabel metal2 s 18906 17325 19014 17435 4 gnd
port 517 nsew
rlabel metal2 s 13434 17895 13542 17971 4 gnd
port 517 nsew
rlabel metal2 s 4698 22855 4806 22965 4 gnd
port 517 nsew
rlabel metal2 s 2202 7625 2310 7701 4 gnd
port 517 nsew
rlabel metal2 s 954 2569 1062 2645 4 gnd
port 517 nsew
rlabel metal2 s 12186 24435 12294 24545 4 gnd
port 517 nsew
rlabel metal2 s 6426 16535 6534 16645 4 gnd
port 517 nsew
rlabel metal2 s 14682 18369 14790 18445 4 gnd
port 517 nsew
rlabel metal2 s 7674 14165 7782 14275 4 gnd
port 517 nsew
rlabel metal2 s 9690 4149 9798 4225 4 gnd
port 517 nsew
rlabel metal2 s 10938 6045 11046 6121 4 gnd
port 517 nsew
rlabel metal2 s 15162 1779 15270 1855 4 gnd
port 517 nsew
rlabel metal2 s 15162 23899 15270 23975 4 gnd
port 517 nsew
rlabel metal2 s 3450 -55 3558 55 4 gnd
port 517 nsew
rlabel metal2 s 18906 16789 19014 16865 4 gnd
port 517 nsew
rlabel metal2 s 13434 19695 13542 19805 4 gnd
port 517 nsew
rlabel metal2 s 9690 11259 9798 11335 4 gnd
port 517 nsew
rlabel metal2 s 17658 1305 17766 1381 4 gnd
port 517 nsew
rlabel metal2 s 4698 14955 4806 15065 4 gnd
port 517 nsew
rlabel metal2 s 18426 16315 18534 16391 4 gnd
port 517 nsew
rlabel metal2 s 10170 16535 10278 16645 4 gnd
port 517 nsew
rlabel metal2 s 19674 5475 19782 5585 4 gnd
port 517 nsew
rlabel metal2 s 10938 18115 11046 18225 4 gnd
port 517 nsew
rlabel metal2 s 2202 5729 2310 5805 4 gnd
port 517 nsew
rlabel metal2 s 19674 16315 19782 16391 4 gnd
port 517 nsew
rlabel metal2 s 2682 17105 2790 17181 4 gnd
port 517 nsew
rlabel metal2 s 13914 13155 14022 13231 4 gnd
port 517 nsew
rlabel metal2 s 16410 7309 16518 7385 4 gnd
port 517 nsew
rlabel metal2 s 954 4939 1062 5015 4 gnd
port 517 nsew
rlabel metal2 s 4698 -55 4806 55 4 gnd
port 517 nsew
rlabel metal2 s 2202 21275 2310 21385 4 gnd
port 517 nsew
rlabel metal2 s 8442 -55 8550 55 4 gnd
port 517 nsew
rlabel metal2 s 14682 23645 14790 23755 4 gnd
port 517 nsew
rlabel metal2 s 17658 199 17766 275 4 gnd
port 517 nsew
rlabel metal2 s 11418 19475 11526 19551 4 gnd
port 517 nsew
rlabel metal2 s 13914 16789 14022 16865 4 gnd
port 517 nsew
rlabel metal2 s 954 10469 1062 10545 4 gnd
port 517 nsew
rlabel metal2 s 5946 18369 6054 18445 4 gnd
port 517 nsew
rlabel metal2 s 15162 22855 15270 22965 4 gnd
port 517 nsew
rlabel metal2 s 13914 515 14022 591 4 gnd
port 517 nsew
rlabel metal2 s 18426 12585 18534 12695 4 gnd
port 517 nsew
rlabel metal2 s 8922 5255 9030 5331 4 gnd
port 517 nsew
rlabel metal2 s 3450 2885 3558 2961 4 gnd
port 517 nsew
rlabel metal2 s 13434 1525 13542 1635 4 gnd
port 517 nsew
rlabel metal2 s 14682 515 14790 591 4 gnd
port 517 nsew
rlabel metal2 s 8442 15525 8550 15601 4 gnd
port 517 nsew
rlabel metal2 s 10938 12049 11046 12125 4 gnd
port 517 nsew
rlabel metal2 s 954 199 1062 275 4 gnd
port 517 nsew
rlabel metal2 s 9690 22635 9798 22711 4 gnd
port 517 nsew
rlabel metal2 s 18426 15209 18534 15285 4 gnd
port 517 nsew
rlabel metal2 s 12186 14955 12294 15065 4 gnd
port 517 nsew
rlabel metal2 s 17658 18685 17766 18761 4 gnd
port 517 nsew
rlabel metal2 s 13434 18905 13542 19015 4 gnd
port 517 nsew
rlabel metal2 s 6426 9425 6534 9535 4 gnd
port 517 nsew
rlabel metal2 s 3450 15745 3558 15855 4 gnd
port 517 nsew
rlabel metal2 s 15162 12049 15270 12125 4 gnd
port 517 nsew
rlabel metal2 s 19674 3895 19782 4005 4 gnd
port 517 nsew
rlabel metal2 s 2202 989 2310 1065 4 gnd
port 517 nsew
rlabel metal2 s 3450 989 3558 1065 4 gnd
port 517 nsew
rlabel metal2 s 10938 1525 11046 1635 4 gnd
port 517 nsew
rlabel metal2 s 13434 11005 13542 11115 4 gnd
port 517 nsew
rlabel metal2 s 15162 23425 15270 23501 4 gnd
port 517 nsew
rlabel metal2 s 186 18369 294 18445 4 gnd
port 517 nsew
rlabel metal2 s 1434 3675 1542 3751 4 gnd
port 517 nsew
rlabel metal2 s 7194 14419 7302 14495 4 gnd
port 517 nsew
rlabel metal2 s 17178 8889 17286 8965 4 gnd
port 517 nsew
rlabel metal2 s 13914 18905 14022 19015 4 gnd
port 517 nsew
rlabel metal2 s 12666 5475 12774 5585 4 gnd
port 517 nsew
rlabel metal2 s 954 22065 1062 22175 4 gnd
port 517 nsew
rlabel metal2 s 2202 10469 2310 10545 4 gnd
port 517 nsew
rlabel metal2 s 4698 24215 4806 24291 4 gnd
port 517 nsew
rlabel metal2 s 5178 12585 5286 12695 4 gnd
port 517 nsew
rlabel metal2 s 13914 9205 14022 9281 4 gnd
port 517 nsew
rlabel metal2 s 8922 6265 9030 6375 4 gnd
port 517 nsew
rlabel metal2 s 1434 989 1542 1065 4 gnd
port 517 nsew
rlabel metal2 s 5946 989 6054 1065 4 gnd
port 517 nsew
rlabel metal2 s 8442 6835 8550 6911 4 gnd
port 517 nsew
rlabel metal2 s 10170 20739 10278 20815 4 gnd
port 517 nsew
rlabel metal2 s 10170 8099 10278 8175 4 gnd
port 517 nsew
rlabel metal2 s 12666 12049 12774 12125 4 gnd
port 517 nsew
rlabel metal2 s 6426 4685 6534 4795 4 gnd
port 517 nsew
rlabel metal2 s 13914 4685 14022 4795 4 gnd
port 517 nsew
rlabel metal2 s 3450 14165 3558 14275 4 gnd
port 517 nsew
rlabel metal2 s 9690 18369 9798 18445 4 gnd
port 517 nsew
rlabel metal2 s 13914 15999 14022 16075 4 gnd
port 517 nsew
rlabel metal2 s 8922 17325 9030 17435 4 gnd
port 517 nsew
rlabel metal2 s 15162 7845 15270 7955 4 gnd
port 517 nsew
rlabel metal2 s 10170 11259 10278 11335 4 gnd
port 517 nsew
rlabel metal2 s 4698 12839 4806 12915 4 gnd
port 517 nsew
rlabel metal2 s 17658 4939 17766 5015 4 gnd
port 517 nsew
rlabel metal2 s 18906 11575 19014 11651 4 gnd
port 517 nsew
rlabel metal2 s 10170 18685 10278 18761 4 gnd
port 517 nsew
rlabel metal2 s 7674 13945 7782 14021 4 gnd
port 517 nsew
rlabel metal2 s 8442 6519 8550 6595 4 gnd
port 517 nsew
rlabel metal2 s 18906 21275 19014 21385 4 gnd
port 517 nsew
rlabel metal2 s 5178 3675 5286 3751 4 gnd
port 517 nsew
rlabel metal2 s 1434 3105 1542 3215 4 gnd
port 517 nsew
rlabel metal2 s 14682 8415 14790 8491 4 gnd
port 517 nsew
rlabel metal2 s 13434 3675 13542 3751 4 gnd
port 517 nsew
rlabel metal2 s 7194 2569 7302 2645 4 gnd
port 517 nsew
rlabel metal2 s 10170 23425 10278 23501 4 gnd
port 517 nsew
rlabel metal2 s 16410 23425 16518 23501 4 gnd
port 517 nsew
rlabel metal2 s 9690 735 9798 845 4 gnd
port 517 nsew
rlabel metal2 s 19674 23899 19782 23975 4 gnd
port 517 nsew
rlabel metal2 s 16410 989 16518 1065 4 gnd
port 517 nsew
rlabel metal2 s 14682 199 14790 275 4 gnd
port 517 nsew
rlabel metal2 s 5178 5729 5286 5805 4 gnd
port 517 nsew
rlabel metal2 s 2682 23899 2790 23975 4 gnd
port 517 nsew
rlabel metal2 s 11418 11259 11526 11335 4 gnd
port 517 nsew
rlabel metal2 s 11418 25225 11526 25335 4 gnd
port 517 nsew
rlabel metal2 s 15162 199 15270 275 4 gnd
port 517 nsew
rlabel metal2 s 13434 8415 13542 8491 4 gnd
port 517 nsew
rlabel metal2 s 13434 16789 13542 16865 4 gnd
port 517 nsew
rlabel metal2 s 10938 19695 11046 19805 4 gnd
port 517 nsew
rlabel metal2 s 8922 17105 9030 17181 4 gnd
port 517 nsew
rlabel metal2 s 2202 24689 2310 24765 4 gnd
port 517 nsew
rlabel metal2 s 7674 10215 7782 10325 4 gnd
port 517 nsew
rlabel metal2 s 18426 25225 18534 25335 4 gnd
port 517 nsew
rlabel metal2 s 13914 2885 14022 2961 4 gnd
port 517 nsew
rlabel metal2 s 18906 3105 19014 3215 4 gnd
port 517 nsew
rlabel metal2 s 13434 -55 13542 55 4 gnd
port 517 nsew
rlabel metal2 s 954 20265 1062 20341 4 gnd
port 517 nsew
rlabel metal2 s 6426 199 6534 275 4 gnd
port 517 nsew
rlabel metal2 s 17178 23899 17286 23975 4 gnd
port 517 nsew
rlabel metal2 s 954 25005 1062 25081 4 gnd
port 517 nsew
rlabel metal2 s 2682 22065 2790 22175 4 gnd
port 517 nsew
rlabel metal2 s 18426 4685 18534 4795 4 gnd
port 517 nsew
rlabel metal2 s 8922 19695 9030 19805 4 gnd
port 517 nsew
rlabel metal2 s 15162 9425 15270 9535 4 gnd
port 517 nsew
rlabel metal2 s 7674 19159 7782 19235 4 gnd
port 517 nsew
rlabel metal2 s 6426 10469 6534 10545 4 gnd
port 517 nsew
rlabel metal2 s 186 14735 294 14811 4 gnd
port 517 nsew
rlabel metal2 s 1434 25005 1542 25081 4 gnd
port 517 nsew
rlabel metal2 s 2682 18905 2790 19015 4 gnd
port 517 nsew
rlabel metal2 s 15930 12365 16038 12441 4 gnd
port 517 nsew
rlabel metal2 s 7194 16789 7302 16865 4 gnd
port 517 nsew
rlabel metal2 s 10170 24435 10278 24545 4 gnd
port 517 nsew
rlabel metal2 s 3450 2569 3558 2645 4 gnd
port 517 nsew
rlabel metal2 s 186 515 294 591 4 gnd
port 517 nsew
rlabel metal2 s 15930 13155 16038 13231 4 gnd
port 517 nsew
rlabel metal2 s 12666 3895 12774 4005 4 gnd
port 517 nsew
rlabel metal2 s 4698 515 4806 591 4 gnd
port 517 nsew
rlabel metal2 s 12666 6519 12774 6595 4 gnd
port 517 nsew
rlabel metal2 s 3450 7625 3558 7701 4 gnd
port 517 nsew
rlabel metal2 s 8922 13375 9030 13485 4 gnd
port 517 nsew
rlabel metal2 s 17658 3675 17766 3751 4 gnd
port 517 nsew
rlabel metal2 s 5946 14955 6054 15065 4 gnd
port 517 nsew
rlabel metal2 s 1434 4465 1542 4541 4 gnd
port 517 nsew
rlabel metal2 s 5946 7055 6054 7165 4 gnd
port 517 nsew
rlabel metal2 s 6426 2315 6534 2425 4 gnd
port 517 nsew
rlabel metal2 s 18906 15209 19014 15285 4 gnd
port 517 nsew
rlabel metal2 s 15162 5255 15270 5331 4 gnd
port 517 nsew
rlabel metal2 s 186 2569 294 2645 4 gnd
port 517 nsew
rlabel metal2 s 16410 12365 16518 12441 4 gnd
port 517 nsew
rlabel metal2 s 17178 22635 17286 22711 4 gnd
port 517 nsew
rlabel metal2 s 3450 8099 3558 8175 4 gnd
port 517 nsew
rlabel metal2 s 2202 21845 2310 21921 4 gnd
port 517 nsew
rlabel metal2 s 2682 9679 2790 9755 4 gnd
port 517 nsew
rlabel metal2 s 11418 6265 11526 6375 4 gnd
port 517 nsew
rlabel metal2 s 4698 3359 4806 3435 4 gnd
port 517 nsew
rlabel metal2 s 186 1305 294 1381 4 gnd
port 517 nsew
rlabel metal2 s 10170 21529 10278 21605 4 gnd
port 517 nsew
rlabel metal2 s 15930 5729 16038 5805 4 gnd
port 517 nsew
rlabel metal2 s 17658 9205 17766 9281 4 gnd
port 517 nsew
rlabel metal2 s 5946 199 6054 275 4 gnd
port 517 nsew
rlabel metal2 s 2202 6045 2310 6121 4 gnd
port 517 nsew
rlabel metal2 s 15162 23645 15270 23755 4 gnd
port 517 nsew
rlabel metal2 s 10170 1525 10278 1635 4 gnd
port 517 nsew
rlabel metal2 s 954 13375 1062 13485 4 gnd
port 517 nsew
rlabel metal2 s 9690 25225 9798 25335 4 gnd
port 517 nsew
rlabel metal2 s 13914 14165 14022 14275 4 gnd
port 517 nsew
rlabel metal2 s 8922 23109 9030 23185 4 gnd
port 517 nsew
rlabel metal2 s 18426 19949 18534 20025 4 gnd
port 517 nsew
rlabel metal2 s 10170 -55 10278 55 4 gnd
port 517 nsew
rlabel metal2 s 15930 2095 16038 2171 4 gnd
port 517 nsew
rlabel metal2 s 5178 15999 5286 16075 4 gnd
port 517 nsew
rlabel metal2 s 186 23109 294 23185 4 gnd
port 517 nsew
rlabel metal2 s 8922 9679 9030 9755 4 gnd
port 517 nsew
rlabel metal2 s 18426 2569 18534 2645 4 gnd
port 517 nsew
rlabel metal2 s 4698 2095 4806 2171 4 gnd
port 517 nsew
rlabel metal2 s 9690 21845 9798 21921 4 gnd
port 517 nsew
rlabel metal2 s 5946 22855 6054 22965 4 gnd
port 517 nsew
rlabel metal2 s 13434 3359 13542 3435 4 gnd
port 517 nsew
rlabel metal2 s 8442 13945 8550 14021 4 gnd
port 517 nsew
rlabel metal2 s 12666 9995 12774 10071 4 gnd
port 517 nsew
rlabel metal2 s 15162 3895 15270 4005 4 gnd
port 517 nsew
rlabel metal2 s 1434 12585 1542 12695 4 gnd
port 517 nsew
rlabel metal2 s 3450 20485 3558 20595 4 gnd
port 517 nsew
rlabel metal2 s 13434 2569 13542 2645 4 gnd
port 517 nsew
rlabel metal2 s 16410 4685 16518 4795 4 gnd
port 517 nsew
rlabel metal2 s 3450 3105 3558 3215 4 gnd
port 517 nsew
rlabel metal2 s 4698 2315 4806 2425 4 gnd
port 517 nsew
rlabel metal2 s 19674 16789 19782 16865 4 gnd
port 517 nsew
rlabel metal2 s 10170 23645 10278 23755 4 gnd
port 517 nsew
rlabel metal2 s 12666 2569 12774 2645 4 gnd
port 517 nsew
rlabel metal2 s 2682 20739 2790 20815 4 gnd
port 517 nsew
rlabel metal2 s 1434 15525 1542 15601 4 gnd
port 517 nsew
rlabel metal2 s 954 24435 1062 24545 4 gnd
port 517 nsew
rlabel metal2 s 5178 199 5286 275 4 gnd
port 517 nsew
rlabel metal2 s 13434 9425 13542 9535 4 gnd
port 517 nsew
rlabel metal2 s 15930 9679 16038 9755 4 gnd
port 517 nsew
rlabel metal2 s 8922 20485 9030 20595 4 gnd
port 517 nsew
rlabel metal2 s 954 9425 1062 9535 4 gnd
port 517 nsew
rlabel metal2 s 1434 5475 1542 5585 4 gnd
port 517 nsew
rlabel metal2 s 9690 7309 9798 7385 4 gnd
port 517 nsew
rlabel metal2 s 11418 15209 11526 15285 4 gnd
port 517 nsew
rlabel metal2 s 14682 989 14790 1065 4 gnd
port 517 nsew
rlabel metal2 s 1434 4685 1542 4795 4 gnd
port 517 nsew
rlabel metal2 s 12186 3895 12294 4005 4 gnd
port 517 nsew
rlabel metal2 s 19674 15525 19782 15601 4 gnd
port 517 nsew
rlabel metal2 s 15162 16315 15270 16391 4 gnd
port 517 nsew
rlabel metal2 s 10938 23899 11046 23975 4 gnd
port 517 nsew
rlabel metal2 s 17178 6835 17286 6911 4 gnd
port 517 nsew
rlabel metal2 s 12186 13945 12294 14021 4 gnd
port 517 nsew
rlabel metal2 s 17178 2885 17286 2961 4 gnd
port 517 nsew
rlabel metal2 s 10938 24215 11046 24291 4 gnd
port 517 nsew
rlabel metal2 s 5178 989 5286 1065 4 gnd
port 517 nsew
rlabel metal2 s 8442 5255 8550 5331 4 gnd
port 517 nsew
rlabel metal2 s 2202 22319 2310 22395 4 gnd
port 517 nsew
rlabel metal2 s 9690 19475 9798 19551 4 gnd
port 517 nsew
rlabel metal2 s 14682 3895 14790 4005 4 gnd
port 517 nsew
rlabel metal2 s 7194 10785 7302 10861 4 gnd
port 517 nsew
rlabel metal2 s 186 15999 294 16075 4 gnd
port 517 nsew
rlabel metal2 s 10170 19159 10278 19235 4 gnd
port 517 nsew
rlabel metal2 s 4698 15525 4806 15601 4 gnd
port 517 nsew
rlabel metal2 s 17658 14955 17766 15065 4 gnd
port 517 nsew
rlabel metal2 s 13914 6265 14022 6375 4 gnd
port 517 nsew
rlabel metal2 s 954 19475 1062 19551 4 gnd
port 517 nsew
rlabel metal2 s 7194 7309 7302 7385 4 gnd
port 517 nsew
rlabel metal2 s 12186 10785 12294 10861 4 gnd
port 517 nsew
rlabel metal2 s 11418 13155 11526 13231 4 gnd
port 517 nsew
rlabel metal2 s 3450 11259 3558 11335 4 gnd
port 517 nsew
rlabel metal2 s 14682 20265 14790 20341 4 gnd
port 517 nsew
rlabel metal2 s 954 15745 1062 15855 4 gnd
port 517 nsew
rlabel metal2 s 10938 14955 11046 15065 4 gnd
port 517 nsew
rlabel metal2 s 14682 12365 14790 12441 4 gnd
port 517 nsew
rlabel metal2 s 18906 13155 19014 13231 4 gnd
port 517 nsew
rlabel metal2 s 17178 1305 17286 1381 4 gnd
port 517 nsew
rlabel metal2 s 186 8635 294 8745 4 gnd
port 517 nsew
rlabel metal2 s 6426 16789 6534 16865 4 gnd
port 517 nsew
rlabel metal2 s 15162 20739 15270 20815 4 gnd
port 517 nsew
rlabel metal2 s 17178 5255 17286 5331 4 gnd
port 517 nsew
rlabel metal2 s 3930 6265 4038 6375 4 gnd
port 517 nsew
rlabel metal2 s 19674 19949 19782 20025 4 gnd
port 517 nsew
rlabel metal2 s 16410 12839 16518 12915 4 gnd
port 517 nsew
rlabel metal2 s 11418 9425 11526 9535 4 gnd
port 517 nsew
rlabel metal2 s 11418 515 11526 591 4 gnd
port 517 nsew
rlabel metal2 s 18426 1525 18534 1635 4 gnd
port 517 nsew
rlabel metal2 s 3930 6835 4038 6911 4 gnd
port 517 nsew
rlabel metal2 s 7674 9425 7782 9535 4 gnd
port 517 nsew
rlabel metal2 s 15930 23109 16038 23185 4 gnd
port 517 nsew
rlabel metal2 s 17178 1779 17286 1855 4 gnd
port 517 nsew
rlabel metal2 s 7674 7055 7782 7165 4 gnd
port 517 nsew
rlabel metal2 s 9690 16789 9798 16865 4 gnd
port 517 nsew
rlabel metal2 s 7674 17579 7782 17655 4 gnd
port 517 nsew
rlabel metal2 s 7194 19949 7302 20025 4 gnd
port 517 nsew
rlabel metal2 s 5178 22319 5286 22395 4 gnd
port 517 nsew
rlabel metal2 s 8442 24215 8550 24291 4 gnd
port 517 nsew
rlabel metal2 s 12186 3105 12294 3215 4 gnd
port 517 nsew
rlabel metal2 s 2202 17895 2310 17971 4 gnd
port 517 nsew
rlabel metal2 s 15930 16315 16038 16391 4 gnd
port 517 nsew
rlabel metal2 s 18906 10469 19014 10545 4 gnd
port 517 nsew
rlabel metal2 s 186 4685 294 4795 4 gnd
port 517 nsew
rlabel metal2 s 19674 25005 19782 25081 4 gnd
port 517 nsew
rlabel metal2 s 7194 199 7302 275 4 gnd
port 517 nsew
rlabel metal2 s 15930 7625 16038 7701 4 gnd
port 517 nsew
rlabel metal2 s 18906 21529 19014 21605 4 gnd
port 517 nsew
rlabel metal2 s 11418 12049 11526 12125 4 gnd
port 517 nsew
rlabel metal2 s 8442 21845 8550 21921 4 gnd
port 517 nsew
rlabel metal2 s 5178 23899 5286 23975 4 gnd
port 517 nsew
rlabel metal2 s 5946 12049 6054 12125 4 gnd
port 517 nsew
rlabel metal2 s 3930 -55 4038 55 4 gnd
port 517 nsew
rlabel metal2 s 8442 10215 8550 10325 4 gnd
port 517 nsew
rlabel metal2 s 13914 -55 14022 55 4 gnd
port 517 nsew
rlabel metal2 s 14682 7625 14790 7701 4 gnd
port 517 nsew
rlabel metal2 s 18906 6519 19014 6595 4 gnd
port 517 nsew
rlabel metal2 s 16410 11575 16518 11651 4 gnd
port 517 nsew
rlabel metal2 s 186 6835 294 6911 4 gnd
port 517 nsew
rlabel metal2 s 17658 10785 17766 10861 4 gnd
port 517 nsew
rlabel metal2 s 13434 6045 13542 6121 4 gnd
port 517 nsew
rlabel metal2 s 1434 10215 1542 10325 4 gnd
port 517 nsew
rlabel metal2 s 16410 22635 16518 22711 4 gnd
port 517 nsew
rlabel metal2 s 14682 14735 14790 14811 4 gnd
port 517 nsew
rlabel metal2 s 18426 13945 18534 14021 4 gnd
port 517 nsew
rlabel metal2 s 19674 5729 19782 5805 4 gnd
port 517 nsew
rlabel metal2 s 3930 3105 4038 3215 4 gnd
port 517 nsew
rlabel metal2 s 8922 23645 9030 23755 4 gnd
port 517 nsew
rlabel metal2 s 3930 7625 4038 7701 4 gnd
port 517 nsew
rlabel metal2 s 9690 21275 9798 21385 4 gnd
port 517 nsew
rlabel metal2 s 12186 19475 12294 19551 4 gnd
port 517 nsew
rlabel metal2 s 11418 10215 11526 10325 4 gnd
port 517 nsew
rlabel metal2 s 10938 13375 11046 13485 4 gnd
port 517 nsew
rlabel metal2 s 10938 14419 11046 14495 4 gnd
port 517 nsew
rlabel metal2 s 2202 20739 2310 20815 4 gnd
port 517 nsew
rlabel metal2 s 1434 12839 1542 12915 4 gnd
port 517 nsew
rlabel metal2 s 2682 8099 2790 8175 4 gnd
port 517 nsew
rlabel metal2 s 13914 4465 14022 4541 4 gnd
port 517 nsew
rlabel metal2 s 13914 25225 14022 25335 4 gnd
port 517 nsew
rlabel metal2 s 15162 18905 15270 19015 4 gnd
port 517 nsew
rlabel metal2 s 17658 11005 17766 11115 4 gnd
port 517 nsew
rlabel metal2 s 7194 6265 7302 6375 4 gnd
port 517 nsew
rlabel metal2 s 18906 5729 19014 5805 4 gnd
port 517 nsew
rlabel metal2 s 6426 24689 6534 24765 4 gnd
port 517 nsew
rlabel metal2 s 7194 7845 7302 7955 4 gnd
port 517 nsew
rlabel metal2 s 4698 2569 4806 2645 4 gnd
port 517 nsew
rlabel metal2 s 8922 8099 9030 8175 4 gnd
port 517 nsew
rlabel metal2 s 7674 19695 7782 19805 4 gnd
port 517 nsew
rlabel metal2 s 2682 4939 2790 5015 4 gnd
port 517 nsew
rlabel metal2 s 17178 2315 17286 2425 4 gnd
port 517 nsew
rlabel metal2 s 10170 2315 10278 2425 4 gnd
port 517 nsew
rlabel metal2 s 4698 23645 4806 23755 4 gnd
port 517 nsew
rlabel metal2 s 8442 15999 8550 16075 4 gnd
port 517 nsew
rlabel metal2 s 8922 12585 9030 12695 4 gnd
port 517 nsew
rlabel metal2 s 18426 12839 18534 12915 4 gnd
port 517 nsew
rlabel metal2 s 9690 9425 9798 9535 4 gnd
port 517 nsew
rlabel metal2 s 10170 8635 10278 8745 4 gnd
port 517 nsew
rlabel metal2 s 3450 9995 3558 10071 4 gnd
port 517 nsew
rlabel metal2 s 2202 21529 2310 21605 4 gnd
port 517 nsew
rlabel metal2 s 954 19949 1062 20025 4 gnd
port 517 nsew
rlabel metal2 s 954 25225 1062 25335 4 gnd
port 517 nsew
rlabel metal2 s 14682 6045 14790 6121 4 gnd
port 517 nsew
rlabel metal2 s 12186 4685 12294 4795 4 gnd
port 517 nsew
rlabel metal2 s 10938 8099 11046 8175 4 gnd
port 517 nsew
rlabel metal2 s 186 23899 294 23975 4 gnd
port 517 nsew
rlabel metal2 s 5946 3105 6054 3215 4 gnd
port 517 nsew
rlabel metal2 s 7674 8099 7782 8175 4 gnd
port 517 nsew
rlabel metal2 s 2682 19475 2790 19551 4 gnd
port 517 nsew
rlabel metal2 s 12666 12839 12774 12915 4 gnd
port 517 nsew
rlabel metal2 s 9690 3675 9798 3751 4 gnd
port 517 nsew
rlabel metal2 s 7194 15745 7302 15855 4 gnd
port 517 nsew
rlabel metal2 s 16410 13629 16518 13705 4 gnd
port 517 nsew
rlabel metal2 s 16410 17895 16518 17971 4 gnd
port 517 nsew
rlabel metal2 s 4698 11795 4806 11905 4 gnd
port 517 nsew
rlabel metal2 s 7194 22635 7302 22711 4 gnd
port 517 nsew
rlabel metal2 s 4698 21529 4806 21605 4 gnd
port 517 nsew
rlabel metal2 s 5946 4939 6054 5015 4 gnd
port 517 nsew
rlabel metal2 s 10170 2569 10278 2645 4 gnd
port 517 nsew
rlabel metal2 s 18906 10785 19014 10861 4 gnd
port 517 nsew
rlabel metal2 s 7194 4465 7302 4541 4 gnd
port 517 nsew
rlabel metal2 s 7194 1525 7302 1635 4 gnd
port 517 nsew
rlabel metal2 s 7674 4939 7782 5015 4 gnd
port 517 nsew
rlabel metal2 s 8442 4149 8550 4225 4 gnd
port 517 nsew
rlabel metal2 s 4698 16315 4806 16391 4 gnd
port 517 nsew
rlabel metal2 s 8442 735 8550 845 4 gnd
port 517 nsew
rlabel metal2 s 1434 16535 1542 16645 4 gnd
port 517 nsew
rlabel metal2 s 1434 14419 1542 14495 4 gnd
port 517 nsew
rlabel metal2 s 5178 21055 5286 21131 4 gnd
port 517 nsew
rlabel metal2 s 2682 5729 2790 5805 4 gnd
port 517 nsew
rlabel metal2 s 6426 19949 6534 20025 4 gnd
port 517 nsew
rlabel metal2 s 7674 21529 7782 21605 4 gnd
port 517 nsew
rlabel metal2 s 16410 7845 16518 7955 4 gnd
port 517 nsew
rlabel metal2 s 954 4465 1062 4541 4 gnd
port 517 nsew
rlabel metal2 s 7674 2095 7782 2171 4 gnd
port 517 nsew
rlabel metal2 s 17178 24435 17286 24545 4 gnd
port 517 nsew
rlabel metal2 s 17658 8889 17766 8965 4 gnd
port 517 nsew
rlabel metal2 s 8922 9425 9030 9535 4 gnd
port 517 nsew
rlabel metal2 s 11418 199 11526 275 4 gnd
port 517 nsew
rlabel metal2 s 15162 21275 15270 21385 4 gnd
port 517 nsew
rlabel metal2 s 19674 12049 19782 12125 4 gnd
port 517 nsew
rlabel metal2 s 19674 4149 19782 4225 4 gnd
port 517 nsew
rlabel metal2 s 4698 7845 4806 7955 4 gnd
port 517 nsew
rlabel metal2 s 17658 24435 17766 24545 4 gnd
port 517 nsew
rlabel metal2 s 13914 20739 14022 20815 4 gnd
port 517 nsew
rlabel metal2 s 10938 21275 11046 21385 4 gnd
port 517 nsew
rlabel metal2 s 954 2315 1062 2425 4 gnd
port 517 nsew
rlabel metal2 s 12666 18115 12774 18225 4 gnd
port 517 nsew
rlabel metal2 s 12666 199 12774 275 4 gnd
port 517 nsew
rlabel metal2 s 9690 13155 9798 13231 4 gnd
port 517 nsew
rlabel metal2 s 12666 19949 12774 20025 4 gnd
port 517 nsew
rlabel metal2 s 3930 12585 4038 12695 4 gnd
port 517 nsew
rlabel metal2 s 10938 2885 11046 2961 4 gnd
port 517 nsew
rlabel metal2 s 8442 12365 8550 12441 4 gnd
port 517 nsew
rlabel metal2 s 15930 14955 16038 15065 4 gnd
port 517 nsew
rlabel metal2 s 7194 12585 7302 12695 4 gnd
port 517 nsew
rlabel metal2 s 5946 14419 6054 14495 4 gnd
port 517 nsew
rlabel metal2 s 14682 22635 14790 22711 4 gnd
port 517 nsew
rlabel metal2 s 6426 21055 6534 21131 4 gnd
port 517 nsew
rlabel metal2 s 7674 10785 7782 10861 4 gnd
port 517 nsew
rlabel metal2 s 186 2885 294 2961 4 gnd
port 517 nsew
rlabel metal2 s 13914 4149 14022 4225 4 gnd
port 517 nsew
rlabel metal2 s 7674 989 7782 1065 4 gnd
port 517 nsew
rlabel metal2 s 5178 4465 5286 4541 4 gnd
port 517 nsew
rlabel metal2 s 4698 199 4806 275 4 gnd
port 517 nsew
rlabel metal2 s 16410 24689 16518 24765 4 gnd
port 517 nsew
rlabel metal2 s 2202 12585 2310 12695 4 gnd
port 517 nsew
rlabel metal2 s 16410 10215 16518 10325 4 gnd
port 517 nsew
rlabel metal2 s 2202 14735 2310 14811 4 gnd
port 517 nsew
rlabel metal2 s 2682 6045 2790 6121 4 gnd
port 517 nsew
rlabel metal2 s 11418 6045 11526 6121 4 gnd
port 517 nsew
rlabel metal2 s 7674 6835 7782 6911 4 gnd
port 517 nsew
rlabel metal2 s 18906 2095 19014 2171 4 gnd
port 517 nsew
rlabel metal2 s 17178 9425 17286 9535 4 gnd
port 517 nsew
rlabel metal2 s 2202 199 2310 275 4 gnd
port 517 nsew
rlabel metal2 s 9690 8099 9798 8175 4 gnd
port 517 nsew
rlabel metal2 s 3930 13945 4038 14021 4 gnd
port 517 nsew
rlabel metal2 s 8922 15525 9030 15601 4 gnd
port 517 nsew
rlabel metal2 s 13914 19159 14022 19235 4 gnd
port 517 nsew
rlabel metal2 s 2202 4939 2310 5015 4 gnd
port 517 nsew
rlabel metal2 s 8922 13155 9030 13231 4 gnd
port 517 nsew
rlabel metal2 s 6426 15209 6534 15285 4 gnd
port 517 nsew
rlabel metal2 s 1434 5255 1542 5331 4 gnd
port 517 nsew
rlabel metal2 s 8922 4465 9030 4541 4 gnd
port 517 nsew
rlabel metal2 s 18906 22635 19014 22711 4 gnd
port 517 nsew
rlabel metal2 s 7194 4939 7302 5015 4 gnd
port 517 nsew
rlabel metal2 s 15930 18115 16038 18225 4 gnd
port 517 nsew
rlabel metal2 s 13434 23425 13542 23501 4 gnd
port 517 nsew
rlabel metal2 s 5178 24689 5286 24765 4 gnd
port 517 nsew
rlabel metal2 s 10170 10215 10278 10325 4 gnd
port 517 nsew
rlabel metal2 s 12666 6265 12774 6375 4 gnd
port 517 nsew
rlabel metal2 s 12666 13155 12774 13231 4 gnd
port 517 nsew
rlabel metal2 s 13434 24689 13542 24765 4 gnd
port 517 nsew
rlabel metal2 s 17178 18905 17286 19015 4 gnd
port 517 nsew
rlabel metal2 s 11418 12365 11526 12441 4 gnd
port 517 nsew
rlabel metal2 s 18426 8415 18534 8491 4 gnd
port 517 nsew
rlabel metal2 s 3450 15209 3558 15285 4 gnd
port 517 nsew
rlabel metal2 s 7674 16315 7782 16391 4 gnd
port 517 nsew
rlabel metal2 s 10938 19949 11046 20025 4 gnd
port 517 nsew
rlabel metal2 s 19674 199 19782 275 4 gnd
port 517 nsew
rlabel metal2 s 16410 2569 16518 2645 4 gnd
port 517 nsew
rlabel metal2 s 16410 8889 16518 8965 4 gnd
port 517 nsew
rlabel metal2 s 10170 9679 10278 9755 4 gnd
port 517 nsew
rlabel metal2 s 7194 20485 7302 20595 4 gnd
port 517 nsew
rlabel metal2 s 9690 6835 9798 6911 4 gnd
port 517 nsew
rlabel metal2 s 3930 11259 4038 11335 4 gnd
port 517 nsew
rlabel metal2 s 14682 23425 14790 23501 4 gnd
port 517 nsew
rlabel metal2 s 8922 12839 9030 12915 4 gnd
port 517 nsew
rlabel metal2 s 15930 22319 16038 22395 4 gnd
port 517 nsew
rlabel metal2 s 7194 14955 7302 15065 4 gnd
port 517 nsew
rlabel metal2 s 8922 6835 9030 6911 4 gnd
port 517 nsew
rlabel metal2 s 6426 9995 6534 10071 4 gnd
port 517 nsew
rlabel metal2 s 11418 25005 11526 25081 4 gnd
port 517 nsew
rlabel metal2 s 10938 25225 11046 25335 4 gnd
port 517 nsew
rlabel metal2 s 10170 13155 10278 13231 4 gnd
port 517 nsew
rlabel metal2 s 18906 6045 19014 6121 4 gnd
port 517 nsew
rlabel metal2 s 13434 23645 13542 23755 4 gnd
port 517 nsew
rlabel metal2 s 6426 5729 6534 5805 4 gnd
port 517 nsew
rlabel metal2 s 4698 10785 4806 10861 4 gnd
port 517 nsew
rlabel metal2 s 6426 13155 6534 13231 4 gnd
port 517 nsew
rlabel metal2 s 18906 24215 19014 24291 4 gnd
port 517 nsew
rlabel metal2 s 18906 1525 19014 1635 4 gnd
port 517 nsew
rlabel metal2 s 4698 1779 4806 1855 4 gnd
port 517 nsew
rlabel metal2 s 15930 18685 16038 18761 4 gnd
port 517 nsew
rlabel metal2 s 12186 12839 12294 12915 4 gnd
port 517 nsew
rlabel metal2 s 7674 8889 7782 8965 4 gnd
port 517 nsew
rlabel metal2 s 954 5729 1062 5805 4 gnd
port 517 nsew
rlabel metal2 s 18426 16535 18534 16645 4 gnd
port 517 nsew
rlabel metal2 s 4698 8635 4806 8745 4 gnd
port 517 nsew
rlabel metal2 s 17658 11575 17766 11651 4 gnd
port 517 nsew
rlabel metal2 s 8442 7625 8550 7701 4 gnd
port 517 nsew
rlabel metal2 s 2682 10469 2790 10545 4 gnd
port 517 nsew
rlabel metal2 s 10170 8415 10278 8491 4 gnd
port 517 nsew
rlabel metal2 s 12186 6265 12294 6375 4 gnd
port 517 nsew
rlabel metal2 s 3450 11795 3558 11905 4 gnd
port 517 nsew
rlabel metal2 s 12186 13155 12294 13231 4 gnd
port 517 nsew
rlabel metal2 s 1434 13375 1542 13485 4 gnd
port 517 nsew
rlabel metal2 s 13914 12365 14022 12441 4 gnd
port 517 nsew
rlabel metal2 s 17178 19695 17286 19805 4 gnd
port 517 nsew
rlabel metal2 s 3450 12585 3558 12695 4 gnd
port 517 nsew
rlabel metal2 s 13914 16315 14022 16391 4 gnd
port 517 nsew
rlabel metal2 s 12186 2095 12294 2171 4 gnd
port 517 nsew
rlabel metal2 s 18426 12049 18534 12125 4 gnd
port 517 nsew
rlabel metal2 s 18426 22319 18534 22395 4 gnd
port 517 nsew
rlabel metal2 s 7674 25005 7782 25081 4 gnd
port 517 nsew
rlabel metal2 s 9690 14735 9798 14811 4 gnd
port 517 nsew
rlabel metal2 s 15162 11575 15270 11651 4 gnd
port 517 nsew
rlabel metal2 s 16410 21275 16518 21385 4 gnd
port 517 nsew
rlabel metal2 s 15930 4149 16038 4225 4 gnd
port 517 nsew
rlabel metal2 s 13434 24435 13542 24545 4 gnd
port 517 nsew
rlabel metal2 s 13914 7625 14022 7701 4 gnd
port 517 nsew
rlabel metal2 s 15162 22065 15270 22175 4 gnd
port 517 nsew
rlabel metal2 s 3450 11005 3558 11115 4 gnd
port 517 nsew
rlabel metal2 s 14682 14165 14790 14275 4 gnd
port 517 nsew
rlabel metal2 s 15162 2885 15270 2961 4 gnd
port 517 nsew
rlabel metal2 s 13914 12049 14022 12125 4 gnd
port 517 nsew
rlabel metal2 s 7194 17325 7302 17435 4 gnd
port 517 nsew
rlabel metal2 s 1434 4939 1542 5015 4 gnd
port 517 nsew
rlabel metal2 s 11418 17105 11526 17181 4 gnd
port 517 nsew
rlabel metal2 s 18426 4939 18534 5015 4 gnd
port 517 nsew
rlabel metal2 s 5946 10469 6054 10545 4 gnd
port 517 nsew
rlabel metal2 s 7194 8635 7302 8745 4 gnd
port 517 nsew
rlabel metal2 s 9690 8415 9798 8491 4 gnd
port 517 nsew
rlabel metal2 s 4698 18369 4806 18445 4 gnd
port 517 nsew
rlabel metal2 s 15930 11005 16038 11115 4 gnd
port 517 nsew
rlabel metal2 s 1434 2569 1542 2645 4 gnd
port 517 nsew
rlabel metal2 s 9690 4465 9798 4541 4 gnd
port 517 nsew
rlabel metal2 s 9690 11575 9798 11651 4 gnd
port 517 nsew
rlabel metal2 s 10938 10785 11046 10861 4 gnd
port 517 nsew
rlabel metal2 s 18426 6265 18534 6375 4 gnd
port 517 nsew
rlabel metal2 s 6426 15525 6534 15601 4 gnd
port 517 nsew
rlabel metal2 s 17658 8099 17766 8175 4 gnd
port 517 nsew
rlabel metal2 s 8442 24689 8550 24765 4 gnd
port 517 nsew
rlabel metal2 s 13434 23899 13542 23975 4 gnd
port 517 nsew
rlabel metal2 s 2682 989 2790 1065 4 gnd
port 517 nsew
rlabel metal2 s 18426 13629 18534 13705 4 gnd
port 517 nsew
rlabel metal2 s 15162 24215 15270 24291 4 gnd
port 517 nsew
rlabel metal2 s 9690 5729 9798 5805 4 gnd
port 517 nsew
rlabel metal2 s 3450 9679 3558 9755 4 gnd
port 517 nsew
rlabel metal2 s 12186 11005 12294 11115 4 gnd
port 517 nsew
rlabel metal2 s 13914 21055 14022 21131 4 gnd
port 517 nsew
rlabel metal2 s 1434 1305 1542 1381 4 gnd
port 517 nsew
rlabel metal2 s 10938 1305 11046 1381 4 gnd
port 517 nsew
rlabel metal2 s 13914 15745 14022 15855 4 gnd
port 517 nsew
rlabel metal2 s 10938 24689 11046 24765 4 gnd
port 517 nsew
rlabel metal2 s 2682 19159 2790 19235 4 gnd
port 517 nsew
rlabel metal2 s 10938 21055 11046 21131 4 gnd
port 517 nsew
rlabel metal2 s 14682 9205 14790 9281 4 gnd
port 517 nsew
rlabel metal2 s 2682 4149 2790 4225 4 gnd
port 517 nsew
rlabel metal2 s 3450 19159 3558 19235 4 gnd
port 517 nsew
rlabel metal2 s 2202 12049 2310 12125 4 gnd
port 517 nsew
rlabel metal2 s 13914 6519 14022 6595 4 gnd
port 517 nsew
rlabel metal2 s 186 14165 294 14275 4 gnd
port 517 nsew
rlabel metal2 s 6426 8415 6534 8491 4 gnd
port 517 nsew
rlabel metal2 s 12186 1525 12294 1635 4 gnd
port 517 nsew
rlabel metal2 s 13914 3105 14022 3215 4 gnd
port 517 nsew
rlabel metal2 s 17178 16789 17286 16865 4 gnd
port 517 nsew
rlabel metal2 s 186 9205 294 9281 4 gnd
port 517 nsew
rlabel metal2 s 17658 21275 17766 21385 4 gnd
port 517 nsew
rlabel metal2 s 12186 25005 12294 25081 4 gnd
port 517 nsew
rlabel metal2 s 18906 3895 19014 4005 4 gnd
port 517 nsew
rlabel metal2 s 10938 5475 11046 5585 4 gnd
port 517 nsew
rlabel metal2 s 186 18905 294 19015 4 gnd
port 517 nsew
rlabel metal2 s 7674 23645 7782 23755 4 gnd
port 517 nsew
rlabel metal2 s 7194 5255 7302 5331 4 gnd
port 517 nsew
rlabel metal2 s 17658 12585 17766 12695 4 gnd
port 517 nsew
rlabel metal2 s 7674 11795 7782 11905 4 gnd
port 517 nsew
rlabel metal2 s 186 19695 294 19805 4 gnd
port 517 nsew
rlabel metal2 s 10938 20739 11046 20815 4 gnd
port 517 nsew
rlabel metal2 s 13914 10215 14022 10325 4 gnd
port 517 nsew
rlabel metal2 s 13434 199 13542 275 4 gnd
port 517 nsew
rlabel metal2 s 19674 4685 19782 4795 4 gnd
port 517 nsew
rlabel metal2 s 3930 9205 4038 9281 4 gnd
port 517 nsew
rlabel metal2 s 5946 24435 6054 24545 4 gnd
port 517 nsew
rlabel metal2 s 2682 13945 2790 14021 4 gnd
port 517 nsew
rlabel metal2 s 954 989 1062 1065 4 gnd
port 517 nsew
rlabel metal2 s 186 15745 294 15855 4 gnd
port 517 nsew
rlabel metal2 s 1434 2315 1542 2425 4 gnd
port 517 nsew
rlabel metal2 s 19674 19159 19782 19235 4 gnd
port 517 nsew
rlabel metal2 s 1434 18905 1542 19015 4 gnd
port 517 nsew
rlabel metal2 s 8442 12049 8550 12125 4 gnd
port 517 nsew
rlabel metal2 s 13914 24689 14022 24765 4 gnd
port 517 nsew
rlabel metal2 s 7194 6835 7302 6911 4 gnd
port 517 nsew
rlabel metal2 s 6426 6265 6534 6375 4 gnd
port 517 nsew
rlabel metal2 s 5946 21055 6054 21131 4 gnd
port 517 nsew
rlabel metal2 s 8442 18115 8550 18225 4 gnd
port 517 nsew
rlabel metal2 s 17178 22319 17286 22395 4 gnd
port 517 nsew
rlabel metal2 s 12666 17325 12774 17435 4 gnd
port 517 nsew
rlabel metal2 s 3450 5475 3558 5585 4 gnd
port 517 nsew
rlabel metal2 s 2682 21275 2790 21385 4 gnd
port 517 nsew
rlabel metal2 s 8442 17895 8550 17971 4 gnd
port 517 nsew
rlabel metal2 s 16410 19695 16518 19805 4 gnd
port 517 nsew
rlabel metal2 s 3450 15999 3558 16075 4 gnd
port 517 nsew
rlabel metal2 s 2682 7309 2790 7385 4 gnd
port 517 nsew
rlabel metal2 s 18426 13155 18534 13231 4 gnd
port 517 nsew
rlabel metal2 s 10938 16315 11046 16391 4 gnd
port 517 nsew
rlabel metal2 s 13434 16535 13542 16645 4 gnd
port 517 nsew
rlabel metal2 s 5946 2315 6054 2425 4 gnd
port 517 nsew
rlabel metal2 s 18426 18685 18534 18761 4 gnd
port 517 nsew
rlabel metal2 s 8922 24215 9030 24291 4 gnd
port 517 nsew
rlabel metal2 s 6426 6519 6534 6595 4 gnd
port 517 nsew
rlabel metal2 s 7674 16789 7782 16865 4 gnd
port 517 nsew
rlabel metal2 s 13914 20265 14022 20341 4 gnd
port 517 nsew
rlabel metal2 s 8442 20485 8550 20595 4 gnd
port 517 nsew
rlabel metal2 s 6426 24435 6534 24545 4 gnd
port 517 nsew
rlabel metal2 s 8442 3895 8550 4005 4 gnd
port 517 nsew
rlabel metal2 s 8922 2569 9030 2645 4 gnd
port 517 nsew
rlabel metal2 s 13914 14735 14022 14811 4 gnd
port 517 nsew
rlabel metal2 s 2682 199 2790 275 4 gnd
port 517 nsew
rlabel metal2 s 8442 4939 8550 5015 4 gnd
port 517 nsew
rlabel metal2 s 8922 16789 9030 16865 4 gnd
port 517 nsew
rlabel metal2 s 7194 16315 7302 16391 4 gnd
port 517 nsew
rlabel metal2 s 5178 10785 5286 10861 4 gnd
port 517 nsew
rlabel metal2 s 8922 18685 9030 18761 4 gnd
port 517 nsew
rlabel metal2 s 11418 5729 11526 5805 4 gnd
port 517 nsew
rlabel metal2 s 15930 13629 16038 13705 4 gnd
port 517 nsew
rlabel metal2 s 3450 11575 3558 11651 4 gnd
port 517 nsew
rlabel metal2 s 1434 25225 1542 25335 4 gnd
port 517 nsew
rlabel metal2 s 2202 13155 2310 13231 4 gnd
port 517 nsew
rlabel metal2 s 7194 17579 7302 17655 4 gnd
port 517 nsew
rlabel metal2 s 186 16789 294 16865 4 gnd
port 517 nsew
rlabel metal2 s 9690 17325 9798 17435 4 gnd
port 517 nsew
rlabel metal2 s 12666 19695 12774 19805 4 gnd
port 517 nsew
rlabel metal2 s 16410 15745 16518 15855 4 gnd
port 517 nsew
rlabel metal2 s 2682 8889 2790 8965 4 gnd
port 517 nsew
rlabel metal2 s 1434 23645 1542 23755 4 gnd
port 517 nsew
rlabel metal2 s 9690 20265 9798 20341 4 gnd
port 517 nsew
rlabel metal2 s 18426 -55 18534 55 4 gnd
port 517 nsew
rlabel metal2 s 954 15999 1062 16075 4 gnd
port 517 nsew
rlabel metal2 s 5178 6835 5286 6911 4 gnd
port 517 nsew
rlabel metal2 s 5946 11259 6054 11335 4 gnd
port 517 nsew
rlabel metal2 s 15162 3675 15270 3751 4 gnd
port 517 nsew
rlabel metal2 s 18426 3675 18534 3751 4 gnd
port 517 nsew
rlabel metal2 s 12666 24689 12774 24765 4 gnd
port 517 nsew
rlabel metal2 s 15162 17895 15270 17971 4 gnd
port 517 nsew
rlabel metal2 s 9690 13945 9798 14021 4 gnd
port 517 nsew
rlabel metal2 s 16410 24215 16518 24291 4 gnd
port 517 nsew
rlabel metal2 s 17658 4465 17766 4541 4 gnd
port 517 nsew
rlabel metal2 s 3450 2315 3558 2425 4 gnd
port 517 nsew
rlabel metal2 s 17658 19159 17766 19235 4 gnd
port 517 nsew
rlabel metal2 s 11418 20739 11526 20815 4 gnd
port 517 nsew
rlabel metal2 s 13434 14735 13542 14811 4 gnd
port 517 nsew
rlabel metal2 s 3450 13629 3558 13705 4 gnd
port 517 nsew
rlabel metal2 s 16410 4465 16518 4541 4 gnd
port 517 nsew
rlabel metal2 s 2682 515 2790 591 4 gnd
port 517 nsew
rlabel metal2 s 5178 7845 5286 7955 4 gnd
port 517 nsew
rlabel metal2 s 15930 16789 16038 16865 4 gnd
port 517 nsew
rlabel metal2 s 19674 5255 19782 5331 4 gnd
port 517 nsew
rlabel metal2 s 12666 13629 12774 13705 4 gnd
port 517 nsew
rlabel metal2 s 16410 4939 16518 5015 4 gnd
port 517 nsew
rlabel metal2 s 7194 2315 7302 2425 4 gnd
port 517 nsew
rlabel metal2 s 10170 21275 10278 21385 4 gnd
port 517 nsew
rlabel metal2 s 12186 11259 12294 11335 4 gnd
port 517 nsew
rlabel metal2 s 2202 11005 2310 11115 4 gnd
port 517 nsew
rlabel metal2 s 8442 2885 8550 2961 4 gnd
port 517 nsew
rlabel metal2 s 16410 3675 16518 3751 4 gnd
port 517 nsew
rlabel metal2 s 5946 18685 6054 18761 4 gnd
port 517 nsew
rlabel metal2 s 13914 6835 14022 6911 4 gnd
port 517 nsew
rlabel metal2 s 18426 23109 18534 23185 4 gnd
port 517 nsew
rlabel metal2 s 12666 11259 12774 11335 4 gnd
port 517 nsew
rlabel metal2 s 13434 20739 13542 20815 4 gnd
port 517 nsew
rlabel metal2 s 2682 17325 2790 17435 4 gnd
port 517 nsew
rlabel metal2 s 7674 14735 7782 14811 4 gnd
port 517 nsew
rlabel metal2 s 4698 6045 4806 6121 4 gnd
port 517 nsew
rlabel metal2 s 8922 1305 9030 1381 4 gnd
port 517 nsew
rlabel metal2 s 12186 19159 12294 19235 4 gnd
port 517 nsew
rlabel metal2 s 5946 7309 6054 7385 4 gnd
port 517 nsew
rlabel metal2 s 4698 25225 4806 25335 4 gnd
port 517 nsew
rlabel metal2 s 18906 4149 19014 4225 4 gnd
port 517 nsew
rlabel metal2 s 15930 735 16038 845 4 gnd
port 517 nsew
rlabel metal2 s 11418 22855 11526 22965 4 gnd
port 517 nsew
rlabel metal2 s 186 3675 294 3751 4 gnd
port 517 nsew
rlabel metal2 s 954 24215 1062 24291 4 gnd
port 517 nsew
rlabel metal2 s 2682 14735 2790 14811 4 gnd
port 517 nsew
rlabel metal2 s 11418 1305 11526 1381 4 gnd
port 517 nsew
rlabel metal2 s 9690 22065 9798 22175 4 gnd
port 517 nsew
rlabel metal2 s 12186 5729 12294 5805 4 gnd
port 517 nsew
rlabel metal2 s 3930 22635 4038 22711 4 gnd
port 517 nsew
rlabel metal2 s 7674 25225 7782 25335 4 gnd
port 517 nsew
rlabel metal2 s 5178 9425 5286 9535 4 gnd
port 517 nsew
rlabel metal2 s 15162 17579 15270 17655 4 gnd
port 517 nsew
rlabel metal2 s 11418 7309 11526 7385 4 gnd
port 517 nsew
rlabel metal2 s 10170 13629 10278 13705 4 gnd
port 517 nsew
rlabel metal2 s 8922 2885 9030 2961 4 gnd
port 517 nsew
rlabel metal2 s 954 17579 1062 17655 4 gnd
port 517 nsew
rlabel metal2 s 5178 19695 5286 19805 4 gnd
port 517 nsew
rlabel metal2 s 8442 24435 8550 24545 4 gnd
port 517 nsew
rlabel metal2 s 12666 10785 12774 10861 4 gnd
port 517 nsew
rlabel metal2 s 3930 9679 4038 9755 4 gnd
port 517 nsew
rlabel metal2 s 12666 15999 12774 16075 4 gnd
port 517 nsew
rlabel metal2 s 2202 18685 2310 18761 4 gnd
port 517 nsew
rlabel metal2 s 5946 7625 6054 7701 4 gnd
port 517 nsew
rlabel metal2 s 10938 7845 11046 7955 4 gnd
port 517 nsew
rlabel metal2 s 2202 4149 2310 4225 4 gnd
port 517 nsew
rlabel metal2 s 15162 8415 15270 8491 4 gnd
port 517 nsew
rlabel metal2 s 8442 21529 8550 21605 4 gnd
port 517 nsew
rlabel metal2 s 15162 19949 15270 20025 4 gnd
port 517 nsew
rlabel metal2 s 2682 1305 2790 1381 4 gnd
port 517 nsew
rlabel metal2 s 14682 21275 14790 21385 4 gnd
port 517 nsew
rlabel metal2 s 1434 515 1542 591 4 gnd
port 517 nsew
rlabel metal2 s 17178 10469 17286 10545 4 gnd
port 517 nsew
rlabel metal2 s 954 7845 1062 7955 4 gnd
port 517 nsew
rlabel metal2 s 2682 13629 2790 13705 4 gnd
port 517 nsew
rlabel metal2 s 8922 7845 9030 7955 4 gnd
port 517 nsew
rlabel metal2 s 13434 3105 13542 3215 4 gnd
port 517 nsew
rlabel metal2 s 2202 515 2310 591 4 gnd
port 517 nsew
rlabel metal2 s 7194 5729 7302 5805 4 gnd
port 517 nsew
rlabel metal2 s 10170 21845 10278 21921 4 gnd
port 517 nsew
rlabel metal2 s 17178 7625 17286 7701 4 gnd
port 517 nsew
rlabel metal2 s 18426 17105 18534 17181 4 gnd
port 517 nsew
rlabel metal2 s 5178 515 5286 591 4 gnd
port 517 nsew
rlabel metal2 s 5946 19695 6054 19805 4 gnd
port 517 nsew
rlabel metal2 s 10938 -55 11046 55 4 gnd
port 517 nsew
rlabel metal2 s 186 25005 294 25081 4 gnd
port 517 nsew
rlabel metal2 s 4698 6265 4806 6375 4 gnd
port 517 nsew
rlabel metal2 s 15930 9995 16038 10071 4 gnd
port 517 nsew
rlabel metal2 s 4698 7625 4806 7701 4 gnd
port 517 nsew
rlabel metal2 s 18906 15525 19014 15601 4 gnd
port 517 nsew
rlabel metal2 s 3450 24435 3558 24545 4 gnd
port 517 nsew
rlabel metal2 s 186 9425 294 9535 4 gnd
port 517 nsew
rlabel metal2 s 7194 7055 7302 7165 4 gnd
port 517 nsew
rlabel metal2 s 8922 14735 9030 14811 4 gnd
port 517 nsew
rlabel metal2 s 4698 21055 4806 21131 4 gnd
port 517 nsew
rlabel metal2 s 4698 11575 4806 11651 4 gnd
port 517 nsew
rlabel metal2 s 15930 12049 16038 12125 4 gnd
port 517 nsew
rlabel metal2 s 17658 14735 17766 14811 4 gnd
port 517 nsew
rlabel metal2 s 5946 14735 6054 14811 4 gnd
port 517 nsew
rlabel metal2 s 9690 16535 9798 16645 4 gnd
port 517 nsew
rlabel metal2 s 12186 5475 12294 5585 4 gnd
port 517 nsew
rlabel metal2 s 7674 3359 7782 3435 4 gnd
port 517 nsew
rlabel metal2 s 19674 13155 19782 13231 4 gnd
port 517 nsew
rlabel metal2 s 10938 9679 11046 9755 4 gnd
port 517 nsew
rlabel metal2 s 8922 23899 9030 23975 4 gnd
port 517 nsew
rlabel metal2 s 13914 19695 14022 19805 4 gnd
port 517 nsew
rlabel metal2 s 2682 14419 2790 14495 4 gnd
port 517 nsew
rlabel metal2 s 5178 8415 5286 8491 4 gnd
port 517 nsew
rlabel metal2 s 9690 23425 9798 23501 4 gnd
port 517 nsew
rlabel metal2 s 17658 22319 17766 22395 4 gnd
port 517 nsew
rlabel metal2 s 12186 17579 12294 17655 4 gnd
port 517 nsew
rlabel metal2 s 3450 14735 3558 14811 4 gnd
port 517 nsew
rlabel metal2 s 5178 15209 5286 15285 4 gnd
port 517 nsew
rlabel metal2 s 5946 8635 6054 8745 4 gnd
port 517 nsew
rlabel metal2 s 6426 3675 6534 3751 4 gnd
port 517 nsew
rlabel metal2 s 7674 6045 7782 6121 4 gnd
port 517 nsew
rlabel metal2 s 5946 13945 6054 14021 4 gnd
port 517 nsew
rlabel metal2 s 12186 7845 12294 7955 4 gnd
port 517 nsew
rlabel metal2 s 5946 3895 6054 4005 4 gnd
port 517 nsew
rlabel metal2 s 8922 15745 9030 15855 4 gnd
port 517 nsew
rlabel metal2 s 12666 9205 12774 9281 4 gnd
port 517 nsew
rlabel metal2 s 18906 15745 19014 15855 4 gnd
port 517 nsew
rlabel metal2 s 17178 21055 17286 21131 4 gnd
port 517 nsew
rlabel metal2 s 186 23645 294 23755 4 gnd
port 517 nsew
rlabel metal2 s 2202 17325 2310 17435 4 gnd
port 517 nsew
rlabel metal2 s 5178 13945 5286 14021 4 gnd
port 517 nsew
rlabel metal2 s 7194 8415 7302 8491 4 gnd
port 517 nsew
rlabel metal2 s 7194 18685 7302 18761 4 gnd
port 517 nsew
rlabel metal2 s 13434 6265 13542 6375 4 gnd
port 517 nsew
rlabel metal2 s 15162 12365 15270 12441 4 gnd
port 517 nsew
rlabel metal2 s 186 16535 294 16645 4 gnd
port 517 nsew
rlabel metal2 s 7194 19695 7302 19805 4 gnd
port 517 nsew
rlabel metal2 s 18426 18369 18534 18445 4 gnd
port 517 nsew
rlabel metal2 s 12186 16789 12294 16865 4 gnd
port 517 nsew
rlabel metal2 s 19674 12839 19782 12915 4 gnd
port 517 nsew
rlabel metal2 s 13434 4465 13542 4541 4 gnd
port 517 nsew
rlabel metal2 s 5178 4939 5286 5015 4 gnd
port 517 nsew
rlabel metal2 s 18906 7845 19014 7955 4 gnd
port 517 nsew
rlabel metal2 s 5178 22855 5286 22965 4 gnd
port 517 nsew
rlabel metal2 s 4698 21845 4806 21921 4 gnd
port 517 nsew
rlabel metal2 s 2682 21529 2790 21605 4 gnd
port 517 nsew
rlabel metal2 s 954 515 1062 591 4 gnd
port 517 nsew
rlabel metal2 s 13434 22635 13542 22711 4 gnd
port 517 nsew
rlabel metal2 s 1434 10785 1542 10861 4 gnd
port 517 nsew
rlabel metal2 s 17178 13629 17286 13705 4 gnd
port 517 nsew
rlabel metal2 s 18426 14735 18534 14811 4 gnd
port 517 nsew
rlabel metal2 s 10170 9205 10278 9281 4 gnd
port 517 nsew
rlabel metal2 s 19674 17895 19782 17971 4 gnd
port 517 nsew
rlabel metal2 s 2682 12365 2790 12441 4 gnd
port 517 nsew
rlabel metal2 s 3930 2885 4038 2961 4 gnd
port 517 nsew
rlabel metal2 s 11418 23899 11526 23975 4 gnd
port 517 nsew
rlabel metal2 s 17658 16789 17766 16865 4 gnd
port 517 nsew
rlabel metal2 s 8922 18115 9030 18225 4 gnd
port 517 nsew
rlabel metal2 s 954 18905 1062 19015 4 gnd
port 517 nsew
rlabel metal2 s 4698 24435 4806 24545 4 gnd
port 517 nsew
rlabel metal2 s 8922 11575 9030 11651 4 gnd
port 517 nsew
rlabel metal2 s 10938 22319 11046 22395 4 gnd
port 517 nsew
rlabel metal2 s 15930 6045 16038 6121 4 gnd
port 517 nsew
rlabel metal2 s 14682 4939 14790 5015 4 gnd
port 517 nsew
rlabel metal2 s 18426 8099 18534 8175 4 gnd
port 517 nsew
rlabel metal2 s 6426 12585 6534 12695 4 gnd
port 517 nsew
rlabel metal2 s 7674 -55 7782 55 4 gnd
port 517 nsew
rlabel metal2 s 5946 21275 6054 21385 4 gnd
port 517 nsew
rlabel metal2 s 10938 8889 11046 8965 4 gnd
port 517 nsew
rlabel metal2 s 15930 11575 16038 11651 4 gnd
port 517 nsew
rlabel metal2 s 954 6265 1062 6375 4 gnd
port 517 nsew
rlabel metal2 s 17658 4685 17766 4795 4 gnd
port 517 nsew
rlabel metal2 s 1434 24435 1542 24545 4 gnd
port 517 nsew
rlabel metal2 s 10170 18369 10278 18445 4 gnd
port 517 nsew
rlabel metal2 s 19674 7055 19782 7165 4 gnd
port 517 nsew
rlabel metal2 s 1434 17895 1542 17971 4 gnd
port 517 nsew
rlabel metal2 s 10938 22635 11046 22711 4 gnd
port 517 nsew
rlabel metal2 s 16410 14165 16518 14275 4 gnd
port 517 nsew
rlabel metal2 s 7674 7845 7782 7955 4 gnd
port 517 nsew
rlabel metal2 s 10938 13629 11046 13705 4 gnd
port 517 nsew
rlabel metal2 s 12186 24215 12294 24291 4 gnd
port 517 nsew
rlabel metal2 s 954 21055 1062 21131 4 gnd
port 517 nsew
rlabel metal2 s 4698 25005 4806 25081 4 gnd
port 517 nsew
rlabel metal2 s 12186 21845 12294 21921 4 gnd
port 517 nsew
rlabel metal2 s 1434 18685 1542 18761 4 gnd
port 517 nsew
rlabel metal2 s 7674 24689 7782 24765 4 gnd
port 517 nsew
<< properties >>
string FIXED_BBOX 0 0 19968 25280
<< end >>
