magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1216 -1260 3724 1750
<< nwell >>
rect 956 0 2464 490
<< pwell >>
rect 411 271 513 462
rect 136 69 788 271
<< scnmos >>
rect 162 155 762 185
<< scpmos >>
rect 1010 155 2410 185
<< ndiff >>
rect 162 237 762 245
rect 162 203 445 237
rect 479 203 762 237
rect 162 185 762 203
rect 162 137 762 155
rect 162 103 445 137
rect 479 103 762 137
rect 162 95 762 103
<< pdiff >>
rect 1010 237 2410 245
rect 1010 203 1693 237
rect 1727 203 2410 237
rect 1010 185 2410 203
rect 1010 137 2410 155
rect 1010 103 1693 137
rect 1727 103 2410 137
rect 1010 95 2410 103
<< ndiffc >>
rect 445 203 479 237
rect 445 103 479 137
<< pdiffc >>
rect 1693 203 1727 237
rect 1693 103 1727 137
<< psubdiff >>
rect 437 412 487 436
rect 437 378 445 412
rect 479 378 487 412
rect 437 354 487 378
<< nsubdiff >>
rect 1685 412 1735 436
rect 1685 378 1693 412
rect 1727 378 1735 412
rect 1685 354 1735 378
<< psubdiffcont >>
rect 445 378 479 412
<< nsubdiffcont >>
rect 1693 378 1727 412
<< poly >>
rect 44 187 110 203
rect 44 153 60 187
rect 94 185 110 187
rect 94 155 162 185
rect 762 155 1010 185
rect 2410 155 2436 185
rect 94 153 110 155
rect 44 137 110 153
<< polycont >>
rect 60 153 94 187
<< locali >>
rect 445 412 479 428
rect 445 362 479 378
rect 1693 412 1727 428
rect 1693 362 1727 378
rect 445 237 479 253
rect 1693 237 1727 253
rect 429 203 445 237
rect 479 203 495 237
rect 1677 203 1693 237
rect 1727 203 1743 237
rect 60 187 94 203
rect 445 187 479 203
rect 1693 187 1727 203
rect 60 137 94 153
rect 429 103 445 137
rect 479 103 1693 137
rect 1727 103 2446 137
<< viali >>
rect 445 378 479 412
rect 1693 378 1727 412
rect 445 203 479 237
rect 1693 203 1727 237
<< metal1 >>
rect 433 412 491 418
rect 433 378 445 412
rect 479 378 491 412
rect 433 372 491 378
rect 1681 412 1739 418
rect 1681 378 1693 412
rect 1727 378 1739 412
rect 1681 372 1739 378
rect 448 243 476 372
rect 1696 243 1724 372
rect 433 237 491 243
rect 433 203 445 237
rect 479 203 491 237
rect 433 197 491 203
rect 1681 237 1739 243
rect 1681 203 1693 237
rect 1727 203 1739 237
rect 1681 197 1739 203
rect 448 0 476 197
rect 1696 0 1724 197
<< labels >>
rlabel locali s 77 170 77 170 4 A
port 2 nsew
rlabel locali s 1437 120 1437 120 4 Z
port 3 nsew
rlabel metal1 s 448 0 476 395 4 gnd
port 5 nsew
rlabel metal1 s 1696 0 1724 395 4 vdd
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2446 41
<< end >>
