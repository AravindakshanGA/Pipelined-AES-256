module s_box_maker (clk, reset, ram_ready, wr_enable, wr_addr, wr_data);
	input clk;
	input reset;
	output reg ram_ready;
	output reg wr_enable;
	output [0:7] wr_addr;
	output [0:7] wr_data;
	
	reg [0:7] count;
	reg [0:7] mem_data_in;
	
	assign wr_addr = count;
	assign wr_data = mem_data_in;
	
	always @(posedge clk) begin
		if(reset == 1'b0) begin
			count <= 8'b0;
			wr_enable <= 1'b0;
			ram_ready <= 1'b0;
		end
		else begin 
			if(count<255) begin 
				wr_enable <= 1'b1;
				ram_ready <= 1'b0;
				if(wr_enable == 1'b1) count <= count + 1'b1;
			end
			else begin
				wr_enable <= 1'b0;
				ram_ready <= 1'b1;
			end
		end
	end

	always @(count) begin
		case (count)
			8'h00: mem_data_in=8'h63;
			8'h01: mem_data_in=8'h7c;
			8'h02: mem_data_in=8'h77;
			8'h03: mem_data_in=8'h7b;
			8'h04: mem_data_in=8'hf2;
			8'h05: mem_data_in=8'h6b;
			8'h06: mem_data_in=8'h6f;
			8'h07: mem_data_in=8'hc5;
			8'h08: mem_data_in=8'h30;
			8'h09: mem_data_in=8'h01;
			8'h0a: mem_data_in=8'h67;
			8'h0b: mem_data_in=8'h2b;
			8'h0c: mem_data_in=8'hfe;
			8'h0d: mem_data_in=8'hd7;
			8'h0e: mem_data_in=8'hab;
			8'h0f: mem_data_in=8'h76;
			8'h10: mem_data_in=8'hca;
			8'h11: mem_data_in=8'h82;
			8'h12: mem_data_in=8'hc9;
			8'h13: mem_data_in=8'h7d;
			8'h14: mem_data_in=8'hfa;
			8'h15: mem_data_in=8'h59;
			8'h16: mem_data_in=8'h47;
			8'h17: mem_data_in=8'hf0;
			8'h18: mem_data_in=8'had;
			8'h19: mem_data_in=8'hd4;
			8'h1a: mem_data_in=8'ha2;
			8'h1b: mem_data_in=8'haf;
			8'h1c: mem_data_in=8'h9c;
			8'h1d: mem_data_in=8'ha4;
			8'h1e: mem_data_in=8'h72;
			8'h1f: mem_data_in=8'hc0;
			8'h20: mem_data_in=8'hb7;
			8'h21: mem_data_in=8'hfd;
			8'h22: mem_data_in=8'h93;
			8'h23: mem_data_in=8'h26;
			8'h24: mem_data_in=8'h36;
			8'h25: mem_data_in=8'h3f;
			8'h26: mem_data_in=8'hf7;
			8'h27: mem_data_in=8'hcc;
			8'h28: mem_data_in=8'h34;
			8'h29: mem_data_in=8'ha5;
			8'h2a: mem_data_in=8'he5;
			8'h2b: mem_data_in=8'hf1;
			8'h2c: mem_data_in=8'h71;
			8'h2d: mem_data_in=8'hd8;
			8'h2e: mem_data_in=8'h31;
			8'h2f: mem_data_in=8'h15;
			8'h30: mem_data_in=8'h04;
			8'h31: mem_data_in=8'hc7;
			8'h32: mem_data_in=8'h23;
			8'h33: mem_data_in=8'hc3;
			8'h34: mem_data_in=8'h18;
			8'h35: mem_data_in=8'h96;
			8'h36: mem_data_in=8'h05;
			8'h37: mem_data_in=8'h9a;
			8'h38: mem_data_in=8'h07;
			8'h39: mem_data_in=8'h12;
			8'h3a: mem_data_in=8'h80;
			8'h3b: mem_data_in=8'he2;
			8'h3c: mem_data_in=8'heb;
			8'h3d: mem_data_in=8'h27;
			8'h3e: mem_data_in=8'hb2;
			8'h3f: mem_data_in=8'h75;
			8'h40: mem_data_in=8'h09;
			8'h41: mem_data_in=8'h83;
			8'h42: mem_data_in=8'h2c;
			8'h43: mem_data_in=8'h1a;
			8'h44: mem_data_in=8'h1b;
			8'h45: mem_data_in=8'h6e;
			8'h46: mem_data_in=8'h5a;
			8'h47: mem_data_in=8'ha0;
			8'h48: mem_data_in=8'h52;
			8'h49: mem_data_in=8'h3b;
			8'h4a: mem_data_in=8'hd6;
			8'h4b: mem_data_in=8'hb3;
			8'h4c: mem_data_in=8'h29;
			8'h4d: mem_data_in=8'he3;
			8'h4e: mem_data_in=8'h2f;
			8'h4f: mem_data_in=8'h84;
			8'h50: mem_data_in=8'h53;
			8'h51: mem_data_in=8'hd1;
			8'h52: mem_data_in=8'h00;
			8'h53: mem_data_in=8'hed;
			8'h54: mem_data_in=8'h20;
			8'h55: mem_data_in=8'hfc;
			8'h56: mem_data_in=8'hb1;
			8'h57: mem_data_in=8'h5b;
			8'h58: mem_data_in=8'h6a;
			8'h59: mem_data_in=8'hcb;
			8'h5a: mem_data_in=8'hbe;
			8'h5b: mem_data_in=8'h39;
			8'h5c: mem_data_in=8'h4a;
			8'h5d: mem_data_in=8'h4c;
			8'h5e: mem_data_in=8'h58;
			8'h5f: mem_data_in=8'hcf;
			8'h60: mem_data_in=8'hd0;
			8'h61: mem_data_in=8'hef;
			8'h62: mem_data_in=8'haa;
			8'h63: mem_data_in=8'hfb;
			8'h64: mem_data_in=8'h43;
			8'h65: mem_data_in=8'h4d;
			8'h66: mem_data_in=8'h33;
			8'h67: mem_data_in=8'h85;
			8'h68: mem_data_in=8'h45;
			8'h69: mem_data_in=8'hf9;
			8'h6a: mem_data_in=8'h02;
			8'h6b: mem_data_in=8'h7f;
			8'h6c: mem_data_in=8'h50;
			8'h6d: mem_data_in=8'h3c;
			8'h6e: mem_data_in=8'h9f;
			8'h6f: mem_data_in=8'ha8;
			8'h70: mem_data_in=8'h51;
			8'h71: mem_data_in=8'ha3;
			8'h72: mem_data_in=8'h40;
			8'h73: mem_data_in=8'h8f;
			8'h74: mem_data_in=8'h92;
			8'h75: mem_data_in=8'h9d;
			8'h76: mem_data_in=8'h38;
			8'h77: mem_data_in=8'hf5;
			8'h78: mem_data_in=8'hbc;
			8'h79: mem_data_in=8'hb6;
			8'h7a: mem_data_in=8'hda;
			8'h7b: mem_data_in=8'h21;
			8'h7c: mem_data_in=8'h10;
			8'h7d: mem_data_in=8'hff;
			8'h7e: mem_data_in=8'hf3;
			8'h7f: mem_data_in=8'hd2;
			8'h80: mem_data_in=8'hcd;
			8'h81: mem_data_in=8'h0c;
			8'h82: mem_data_in=8'h13;
			8'h83: mem_data_in=8'hec;
			8'h84: mem_data_in=8'h5f;
			8'h85: mem_data_in=8'h97;
			8'h86: mem_data_in=8'h44;
			8'h87: mem_data_in=8'h17;
			8'h88: mem_data_in=8'hc4;
			8'h89: mem_data_in=8'ha7;
			8'h8a: mem_data_in=8'h7e;
			8'h8b: mem_data_in=8'h3d;
			8'h8c: mem_data_in=8'h64;
			8'h8d: mem_data_in=8'h5d;
			8'h8e: mem_data_in=8'h19;
			8'h8f: mem_data_in=8'h73;
			8'h90: mem_data_in=8'h60;
			8'h91: mem_data_in=8'h81;
			8'h92: mem_data_in=8'h4f;
			8'h93: mem_data_in=8'hdc;
			8'h94: mem_data_in=8'h22;
			8'h95: mem_data_in=8'h2a;
			8'h96: mem_data_in=8'h90;
			8'h97: mem_data_in=8'h88;
			8'h98: mem_data_in=8'h46;
			8'h99: mem_data_in=8'hee;
			8'h9a: mem_data_in=8'hb8;
			8'h9b: mem_data_in=8'h14;
			8'h9c: mem_data_in=8'hde;
			8'h9d: mem_data_in=8'h5e;
			8'h9e: mem_data_in=8'h0b;
			8'h9f: mem_data_in=8'hdb;
			8'ha0: mem_data_in=8'he0;
			8'ha1: mem_data_in=8'h32;
			8'ha2: mem_data_in=8'h3a;
			8'ha3: mem_data_in=8'h0a;
			8'ha4: mem_data_in=8'h49;
			8'ha5: mem_data_in=8'h06;
			8'ha6: mem_data_in=8'h24;
			8'ha7: mem_data_in=8'h5c;
			8'ha8: mem_data_in=8'hc2;
			8'ha9: mem_data_in=8'hd3;
			8'haa: mem_data_in=8'hac;
			8'hab: mem_data_in=8'h62;
			8'hac: mem_data_in=8'h91;
			8'had: mem_data_in=8'h95;
			8'hae: mem_data_in=8'he4;
			8'haf: mem_data_in=8'h79;
			8'hb0: mem_data_in=8'he7;
			8'hb1: mem_data_in=8'hc8;
			8'hb2: mem_data_in=8'h37;
			8'hb3: mem_data_in=8'h6d;
			8'hb4: mem_data_in=8'h8d;
			8'hb5: mem_data_in=8'hd5;
			8'hb6: mem_data_in=8'h4e;
			8'hb7: mem_data_in=8'ha9;
			8'hb8: mem_data_in=8'h6c;
			8'hb9: mem_data_in=8'h56;
			8'hba: mem_data_in=8'hf4;
			8'hbb: mem_data_in=8'hea;
			8'hbc: mem_data_in=8'h65;
			8'hbd: mem_data_in=8'h7a;
			8'hbe: mem_data_in=8'hae;
			8'hbf: mem_data_in=8'h08;
			8'hc0: mem_data_in=8'hba;
			8'hc1: mem_data_in=8'h78;
			8'hc2: mem_data_in=8'h25;
			8'hc3: mem_data_in=8'h2e;
			8'hc4: mem_data_in=8'h1c;
			8'hc5: mem_data_in=8'ha6;
			8'hc6: mem_data_in=8'hb4;
			8'hc7: mem_data_in=8'hc6;
			8'hc8: mem_data_in=8'he8;
			8'hc9: mem_data_in=8'hdd;
			8'hca: mem_data_in=8'h74;
			8'hcb: mem_data_in=8'h1f;
			8'hcc: mem_data_in=8'h4b;
			8'hcd: mem_data_in=8'hbd;
			8'hce: mem_data_in=8'h8b;
			8'hcf: mem_data_in=8'h8a;
			8'hd0: mem_data_in=8'h70;
			8'hd1: mem_data_in=8'h3e;
			8'hd2: mem_data_in=8'hb5;
			8'hd3: mem_data_in=8'h66;
			8'hd4: mem_data_in=8'h48;
			8'hd5: mem_data_in=8'h03;
			8'hd6: mem_data_in=8'hf6;
			8'hd7: mem_data_in=8'h0e;
			8'hd8: mem_data_in=8'h61;
			8'hd9: mem_data_in=8'h35;
			8'hda: mem_data_in=8'h57;
			8'hdb: mem_data_in=8'hb9;
			8'hdc: mem_data_in=8'h86;
			8'hdd: mem_data_in=8'hc1;
			8'hde: mem_data_in=8'h1d;
			8'hdf: mem_data_in=8'h9e;
			8'he0: mem_data_in=8'he1;
			8'he1: mem_data_in=8'hf8;
			8'he2: mem_data_in=8'h98;
			8'he3: mem_data_in=8'h11;
			8'he4: mem_data_in=8'h69;
			8'he5: mem_data_in=8'hd9;
			8'he6: mem_data_in=8'h8e;
			8'he7: mem_data_in=8'h94;
			8'he8: mem_data_in=8'h9b;
			8'he9: mem_data_in=8'h1e;
			8'hea: mem_data_in=8'h87;
			8'heb: mem_data_in=8'he9;
			8'hec: mem_data_in=8'hce;
			8'hed: mem_data_in=8'h55;
			8'hee: mem_data_in=8'h28;
			8'hef: mem_data_in=8'hdf;
			8'hf0: mem_data_in=8'h8c;
			8'hf1: mem_data_in=8'ha1;
			8'hf2: mem_data_in=8'h89;
			8'hf3: mem_data_in=8'h0d;
			8'hf4: mem_data_in=8'hbf;
			8'hf5: mem_data_in=8'he6;
			8'hf6: mem_data_in=8'h42;
			8'hf7: mem_data_in=8'h68;
			8'hf8: mem_data_in=8'h41;
			8'hf9: mem_data_in=8'h99;
			8'hfa: mem_data_in=8'h2d;
			8'hfb: mem_data_in=8'h0f;
			8'hfc: mem_data_in=8'hb0;
			8'hfd: mem_data_in=8'h54;
			8'hfe: mem_data_in=8'hbb;
			8'hff: mem_data_in=8'h16;
		endcase
	end
endmodule