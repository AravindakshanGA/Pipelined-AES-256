magic
tech sky130A
magscale 1 2
timestamp 1543373569
<< checkpaint >>
rect -1260 -1750 11949 26605
<< locali >>
rect 6844 25143 7045 25177
rect 10643 25143 10677 25177
rect 7011 24998 7045 25143
rect 7011 24964 7436 24998
rect 7011 24772 7436 24806
rect 7011 24627 7045 24772
rect 6844 24593 7045 24627
rect 10643 24593 10677 24627
rect 6844 24353 7045 24387
rect 10643 24353 10677 24387
rect 7011 24208 7045 24353
rect 7011 24174 7436 24208
rect 7011 23982 7436 24016
rect 7011 23837 7045 23982
rect 6844 23803 7045 23837
rect 10643 23803 10677 23837
rect 6844 23563 7045 23597
rect 10643 23563 10677 23597
rect 7011 23418 7045 23563
rect 7011 23384 7436 23418
rect 7011 23192 7436 23226
rect 7011 23047 7045 23192
rect 6844 23013 7045 23047
rect 10643 23013 10677 23047
rect 6844 22773 7045 22807
rect 10643 22773 10677 22807
rect 7011 22628 7045 22773
rect 7011 22594 7436 22628
rect 7011 22402 7436 22436
rect 7011 22257 7045 22402
rect 6844 22223 7045 22257
rect 10643 22223 10677 22257
rect 6844 21983 7045 22017
rect 10643 21983 10677 22017
rect 7011 21838 7045 21983
rect 7011 21804 7436 21838
rect 7011 21612 7436 21646
rect 7011 21467 7045 21612
rect 6844 21433 7045 21467
rect 10643 21433 10677 21467
rect 6844 21193 7045 21227
rect 10643 21193 10677 21227
rect 7011 21048 7045 21193
rect 7011 21014 7436 21048
rect 7011 20822 7436 20856
rect 7011 20677 7045 20822
rect 6844 20643 7045 20677
rect 10643 20643 10677 20677
rect 6844 20403 7045 20437
rect 10643 20403 10677 20437
rect 7011 20258 7045 20403
rect 7011 20224 7436 20258
rect 7011 20032 7436 20066
rect 7011 19887 7045 20032
rect 6844 19853 7045 19887
rect 10643 19853 10677 19887
rect 6844 19613 7045 19647
rect 10643 19613 10677 19647
rect 7011 19468 7045 19613
rect 7011 19434 7436 19468
rect 7011 19242 7436 19276
rect 7011 19097 7045 19242
rect 6844 19063 7045 19097
rect 10643 19063 10677 19097
rect 6844 18823 7045 18857
rect 10643 18823 10677 18857
rect 7011 18678 7045 18823
rect 7011 18644 7436 18678
rect 7011 18452 7436 18486
rect 7011 18307 7045 18452
rect 6844 18273 7045 18307
rect 10643 18273 10677 18307
rect 6844 18033 7045 18067
rect 10643 18033 10677 18067
rect 7011 17888 7045 18033
rect 7011 17854 7436 17888
rect 7011 17662 7436 17696
rect 7011 17517 7045 17662
rect 6844 17483 7045 17517
rect 10643 17483 10677 17517
rect 6844 17243 7045 17277
rect 10643 17243 10677 17277
rect 7011 17098 7045 17243
rect 7011 17064 7436 17098
rect 7011 16872 7436 16906
rect 7011 16727 7045 16872
rect 6844 16693 7045 16727
rect 10643 16693 10677 16727
rect 6844 16453 7045 16487
rect 10643 16453 10677 16487
rect 7011 16308 7045 16453
rect 7011 16274 7436 16308
rect 7011 16082 7436 16116
rect 7011 15937 7045 16082
rect 6844 15903 7045 15937
rect 10643 15903 10677 15937
rect 6844 15663 7045 15697
rect 10643 15663 10677 15697
rect 7011 15518 7045 15663
rect 7011 15484 7436 15518
rect 7011 15292 7436 15326
rect 7011 15147 7045 15292
rect 6844 15113 7045 15147
rect 10643 15113 10677 15147
rect 6844 14873 7045 14907
rect 10643 14873 10677 14907
rect 7011 14728 7045 14873
rect 7011 14694 7436 14728
rect 7011 14502 7436 14536
rect 7011 14357 7045 14502
rect 6844 14323 7045 14357
rect 10643 14323 10677 14357
rect 6844 14083 7045 14117
rect 10643 14083 10677 14117
rect 7011 13938 7045 14083
rect 7011 13904 7436 13938
rect 7011 13712 7436 13746
rect 7011 13567 7045 13712
rect 6844 13533 7045 13567
rect 10643 13533 10677 13567
rect 6844 13293 7045 13327
rect 10643 13293 10677 13327
rect 7011 13148 7045 13293
rect 7011 13114 7436 13148
rect 7011 12922 7436 12956
rect 7011 12777 7045 12922
rect 6844 12743 7045 12777
rect 10643 12743 10677 12777
rect 6844 12503 7045 12537
rect 10643 12503 10677 12537
rect 7011 12358 7045 12503
rect 7011 12324 7436 12358
rect 7011 12132 7436 12166
rect 7011 11987 7045 12132
rect 6844 11953 7045 11987
rect 10643 11953 10677 11987
rect 6844 11713 7045 11747
rect 10643 11713 10677 11747
rect 7011 11568 7045 11713
rect 7011 11534 7436 11568
rect 7011 11342 7436 11376
rect 7011 11197 7045 11342
rect 6844 11163 7045 11197
rect 10643 11163 10677 11197
rect 6844 10923 7045 10957
rect 10643 10923 10677 10957
rect 7011 10778 7045 10923
rect 7011 10744 7436 10778
rect 7011 10552 7436 10586
rect 7011 10407 7045 10552
rect 6844 10373 7045 10407
rect 10643 10373 10677 10407
rect 6844 10133 7045 10167
rect 10643 10133 10677 10167
rect 7011 9988 7045 10133
rect 7011 9954 7436 9988
rect 7011 9762 7436 9796
rect 7011 9617 7045 9762
rect 6844 9583 7045 9617
rect 10643 9583 10677 9617
rect 6844 9343 7045 9377
rect 10643 9343 10677 9377
rect 7011 9198 7045 9343
rect 7011 9164 7436 9198
rect 7011 8972 7436 9006
rect 7011 8827 7045 8972
rect 6844 8793 7045 8827
rect 10643 8793 10677 8827
rect 6844 8553 7045 8587
rect 10643 8553 10677 8587
rect 7011 8408 7045 8553
rect 7011 8374 7436 8408
rect 7011 8182 7436 8216
rect 7011 8037 7045 8182
rect 6844 8003 7045 8037
rect 10643 8003 10677 8037
rect 6844 7763 7045 7797
rect 10643 7763 10677 7797
rect 7011 7618 7045 7763
rect 7011 7584 7436 7618
rect 7011 7392 7436 7426
rect 7011 7247 7045 7392
rect 6844 7213 7045 7247
rect 10643 7213 10677 7247
rect 6844 6973 7045 7007
rect 10643 6973 10677 7007
rect 7011 6828 7045 6973
rect 7011 6794 7436 6828
rect 7011 6602 7436 6636
rect 7011 6457 7045 6602
rect 6844 6423 7045 6457
rect 10643 6423 10677 6457
rect 6844 6183 7045 6217
rect 10643 6183 10677 6217
rect 7011 6038 7045 6183
rect 7011 6004 7436 6038
rect 7011 5812 7436 5846
rect 7011 5667 7045 5812
rect 6844 5633 7045 5667
rect 10643 5633 10677 5667
rect 6844 5393 7045 5427
rect 10643 5393 10677 5427
rect 7011 5248 7045 5393
rect 7011 5214 7436 5248
rect 7011 5022 7436 5056
rect 7011 4877 7045 5022
rect 6844 4843 7045 4877
rect 10643 4843 10677 4877
rect 6844 4603 7045 4637
rect 10643 4603 10677 4637
rect 7011 4458 7045 4603
rect 7011 4424 7436 4458
rect 7011 4232 7436 4266
rect 7011 4087 7045 4232
rect 6844 4053 7045 4087
rect 10643 4053 10677 4087
rect 6844 3813 7045 3847
rect 10643 3813 10677 3847
rect 7011 3668 7045 3813
rect 7011 3634 7436 3668
rect 7011 3442 7436 3476
rect 7011 3297 7045 3442
rect 6844 3263 7045 3297
rect 10643 3263 10677 3297
rect 6844 3023 7045 3057
rect 10643 3023 10677 3057
rect 7011 2878 7045 3023
rect 7011 2844 7436 2878
rect 7011 2652 7436 2686
rect 7011 2507 7045 2652
rect 6844 2473 7045 2507
rect 10643 2473 10677 2507
rect 6844 2233 7045 2267
rect 10643 2233 10677 2267
rect 7011 2088 7045 2233
rect 7011 2054 7436 2088
rect 7011 1862 7436 1896
rect 7011 1717 7045 1862
rect 6844 1683 7045 1717
rect 10643 1683 10677 1717
rect 6844 1443 7045 1477
rect 10643 1443 10677 1477
rect 7011 1298 7045 1443
rect 7011 1264 7436 1298
rect 7011 1072 7436 1106
rect 7011 927 7045 1072
rect 6844 893 7045 927
rect 10643 893 10677 927
rect 6844 653 7045 687
rect 10643 653 10677 687
rect 7011 508 7045 653
rect 7011 474 7436 508
rect 7011 282 7436 316
rect 7011 137 7045 282
rect 6844 103 7045 137
rect 10643 103 10677 137
rect 8654 -137 10671 -103
rect 7195 -174 7229 -158
rect 7229 -208 7452 -174
rect 7195 -224 7229 -208
rect 7435 -282 7469 -266
rect 7435 -332 7469 -316
<< viali >>
rect 7195 -208 7229 -174
rect 7435 -316 7469 -282
<< metal1 >>
rect 19 0 47 6320
rect 99 0 127 6320
rect 179 0 207 6320
rect 259 0 287 6320
rect 339 0 367 6320
rect 419 0 447 6320
rect 7180 -217 7186 -165
rect 7238 -217 7244 -165
rect 7420 -325 7426 -273
rect 7478 -325 7484 -273
rect 8019 -402 8069 32
rect 9921 -395 9949 0
<< via1 >>
rect 7186 -174 7238 -165
rect 7186 -208 7195 -174
rect 7195 -208 7229 -174
rect 7229 -208 7238 -174
rect 7186 -217 7238 -208
rect 7426 -282 7478 -273
rect 7426 -316 7435 -282
rect 7435 -316 7469 -282
rect 7469 -316 7478 -282
rect 7426 -325 7478 -316
<< metal2 >>
rect 7184 -163 7240 -154
rect 7184 -228 7240 -219
rect 7438 -267 7466 0
rect 7426 -273 7478 -267
rect 7426 -331 7478 -325
<< via2 >>
rect 7184 -165 7240 -163
rect 7184 -217 7186 -165
rect 7186 -217 7238 -165
rect 7238 -217 7240 -165
rect 7184 -219 7240 -217
<< metal3 >>
rect 2290 5883 2388 5981
rect 2715 5883 2813 5981
rect 3094 5876 3192 5974
rect 3490 5876 3588 5974
rect 996 5086 1094 5184
rect 1392 5086 1490 5184
rect 2290 5093 2388 5191
rect 2715 5093 2813 5191
rect 3094 5086 3192 5184
rect 3490 5086 3588 5184
rect 2290 3513 2388 3611
rect 2715 3513 2813 3611
rect 3094 3506 3192 3604
rect 3490 3506 3588 3604
rect 996 2716 1094 2814
rect 1392 2716 1490 2814
rect 2290 2723 2388 2821
rect 2715 2723 2813 2821
rect 3094 2716 3192 2814
rect 3490 2716 3588 2814
rect 2290 1143 2388 1241
rect 2715 1143 2813 1241
rect 3094 1136 3192 1234
rect 3490 1136 3588 1234
rect 996 346 1094 444
rect 1392 346 1490 444
rect 2290 353 2388 451
rect 2715 353 2813 451
rect 3094 346 3192 444
rect 3490 346 3588 444
rect 7163 -163 7261 -142
rect 7163 -219 7184 -163
rect 7240 -219 7261 -163
rect 7163 -240 7261 -219
<< metal4 >>
rect 5022 -33 5088 25341
rect 5494 -33 5560 25341
rect 5926 -33 5992 25341
rect 6270 -33 6336 25341
rect 6694 -33 6760 25341
rect 7586 -63 7652 25343
rect 8011 -65 8077 25345
rect 8654 -33 8720 25313
rect 9902 -33 9968 25313
use subbyte2_and2_dec_0  subbyte2_and2_dec_0_0
timestamp 1543373570
transform 1 0 7349 0 -1 0
box 70 -56 3340 490
use subbyte2_hierarchical_decoder  subbyte2_hierarchical_decoder_0
timestamp 1543373569
transform 1 0 0 0 1 0
box 0 -60 6879 25341
use subbyte2_wordline_driver_array  subbyte2_wordline_driver_array_0
timestamp 1543373570
transform 1 0 6861 0 1 0
box 558 -65 3828 25345
<< labels >>
rlabel metal1 s 19 0 47 6320 4 addr_0
port 3 nsew
rlabel metal1 s 99 0 127 6320 4 addr_1
port 5 nsew
rlabel metal1 s 179 0 207 6320 4 addr_2
port 7 nsew
rlabel metal1 s 259 0 287 6320 4 addr_3
port 9 nsew
rlabel metal1 s 339 0 367 6320 4 addr_4
port 11 nsew
rlabel metal1 s 419 0 447 6320 4 addr_5
port 13 nsew
rlabel locali s 10660 120 10660 120 4 wl_0
port 14 nsew
rlabel locali s 10660 670 10660 670 4 wl_1
port 15 nsew
rlabel locali s 10660 910 10660 910 4 wl_2
port 16 nsew
rlabel locali s 10660 1460 10660 1460 4 wl_3
port 17 nsew
rlabel locali s 10660 1700 10660 1700 4 wl_4
port 18 nsew
rlabel locali s 10660 2250 10660 2250 4 wl_5
port 19 nsew
rlabel locali s 10660 2490 10660 2490 4 wl_6
port 20 nsew
rlabel locali s 10660 3040 10660 3040 4 wl_7
port 21 nsew
rlabel locali s 10660 3280 10660 3280 4 wl_8
port 22 nsew
rlabel locali s 10660 3830 10660 3830 4 wl_9
port 23 nsew
rlabel locali s 10660 4070 10660 4070 4 wl_10
port 24 nsew
rlabel locali s 10660 4620 10660 4620 4 wl_11
port 25 nsew
rlabel locali s 10660 4860 10660 4860 4 wl_12
port 26 nsew
rlabel locali s 10660 5410 10660 5410 4 wl_13
port 27 nsew
rlabel locali s 10660 5650 10660 5650 4 wl_14
port 28 nsew
rlabel locali s 10660 6200 10660 6200 4 wl_15
port 29 nsew
rlabel locali s 10660 6440 10660 6440 4 wl_16
port 30 nsew
rlabel locali s 10660 6990 10660 6990 4 wl_17
port 31 nsew
rlabel locali s 10660 7230 10660 7230 4 wl_18
port 32 nsew
rlabel locali s 10660 7780 10660 7780 4 wl_19
port 33 nsew
rlabel locali s 10660 8020 10660 8020 4 wl_20
port 34 nsew
rlabel locali s 10660 8570 10660 8570 4 wl_21
port 35 nsew
rlabel locali s 10660 8810 10660 8810 4 wl_22
port 36 nsew
rlabel locali s 10660 9360 10660 9360 4 wl_23
port 37 nsew
rlabel locali s 10660 9600 10660 9600 4 wl_24
port 38 nsew
rlabel locali s 10660 10150 10660 10150 4 wl_25
port 39 nsew
rlabel locali s 10660 10390 10660 10390 4 wl_26
port 40 nsew
rlabel locali s 10660 10940 10660 10940 4 wl_27
port 41 nsew
rlabel locali s 10660 11180 10660 11180 4 wl_28
port 42 nsew
rlabel locali s 10660 11730 10660 11730 4 wl_29
port 43 nsew
rlabel locali s 10660 11970 10660 11970 4 wl_30
port 44 nsew
rlabel locali s 10660 12520 10660 12520 4 wl_31
port 45 nsew
rlabel locali s 10660 12760 10660 12760 4 wl_32
port 46 nsew
rlabel locali s 10660 13310 10660 13310 4 wl_33
port 47 nsew
rlabel locali s 10660 13550 10660 13550 4 wl_34
port 48 nsew
rlabel locali s 10660 14100 10660 14100 4 wl_35
port 49 nsew
rlabel locali s 10660 14340 10660 14340 4 wl_36
port 50 nsew
rlabel locali s 10660 14890 10660 14890 4 wl_37
port 51 nsew
rlabel locali s 10660 15130 10660 15130 4 wl_38
port 52 nsew
rlabel locali s 10660 15680 10660 15680 4 wl_39
port 53 nsew
rlabel locali s 10660 15920 10660 15920 4 wl_40
port 54 nsew
rlabel locali s 10660 16470 10660 16470 4 wl_41
port 55 nsew
rlabel locali s 10660 16710 10660 16710 4 wl_42
port 56 nsew
rlabel locali s 10660 17260 10660 17260 4 wl_43
port 57 nsew
rlabel locali s 10660 17500 10660 17500 4 wl_44
port 58 nsew
rlabel locali s 10660 18050 10660 18050 4 wl_45
port 59 nsew
rlabel locali s 10660 18290 10660 18290 4 wl_46
port 60 nsew
rlabel locali s 10660 18840 10660 18840 4 wl_47
port 61 nsew
rlabel locali s 10660 19080 10660 19080 4 wl_48
port 62 nsew
rlabel locali s 10660 19630 10660 19630 4 wl_49
port 63 nsew
rlabel locali s 10660 19870 10660 19870 4 wl_50
port 64 nsew
rlabel locali s 10660 20420 10660 20420 4 wl_51
port 65 nsew
rlabel locali s 10660 20660 10660 20660 4 wl_52
port 66 nsew
rlabel locali s 10660 21210 10660 21210 4 wl_53
port 67 nsew
rlabel locali s 10660 21450 10660 21450 4 wl_54
port 68 nsew
rlabel locali s 10660 22000 10660 22000 4 wl_55
port 69 nsew
rlabel locali s 10660 22240 10660 22240 4 wl_56
port 70 nsew
rlabel locali s 10660 22790 10660 22790 4 wl_57
port 71 nsew
rlabel locali s 10660 23030 10660 23030 4 wl_58
port 72 nsew
rlabel locali s 10660 23580 10660 23580 4 wl_59
port 73 nsew
rlabel locali s 10660 23820 10660 23820 4 wl_60
port 74 nsew
rlabel locali s 10660 24370 10660 24370 4 wl_61
port 75 nsew
rlabel locali s 10660 24610 10660 24610 4 wl_62
port 76 nsew
rlabel locali s 10660 25160 10660 25160 4 wl_63
port 77 nsew
rlabel locali s 9662 -120 9662 -120 4 rbl_wl
port 78 nsew
rlabel metal2 s 7438 -313 7466 -285 4 wl_en
port 80 nsew
rlabel metal3 s 3490 1136 3588 1234 4 vdd
port 82 nsew
rlabel metal3 s 2715 5093 2813 5191 4 vdd
port 82 nsew
rlabel metal3 s 2715 1143 2813 1241 4 vdd
port 82 nsew
rlabel metal3 s 1392 346 1490 444 4 vdd
port 82 nsew
rlabel metal3 s 1392 5086 1490 5184 4 vdd
port 82 nsew
rlabel metal3 s 3490 2716 3588 2814 4 vdd
port 82 nsew
rlabel metal3 s 2715 2723 2813 2821 4 vdd
port 82 nsew
rlabel metal4 s 8011 -65 8077 25345 4 vdd
port 82 nsew
rlabel metal3 s 3490 5876 3588 5974 4 vdd
port 82 nsew
rlabel metal3 s 3490 5086 3588 5184 4 vdd
port 82 nsew
rlabel metal3 s 3490 3506 3588 3604 4 vdd
port 82 nsew
rlabel metal3 s 7163 -240 7261 -142 4 vdd
port 82 nsew
rlabel metal1 s 9921 -395 9949 0 4 vdd
port 82 nsew
rlabel metal3 s 2715 5883 2813 5981 4 vdd
port 82 nsew
rlabel metal1 s 8019 -402 8069 32 4 vdd
port 82 nsew
rlabel metal3 s 3490 346 3588 444 4 vdd
port 82 nsew
rlabel metal4 s 6694 -33 6760 25341 4 vdd
port 82 nsew
rlabel metal4 s 5494 -33 5560 25341 4 vdd
port 82 nsew
rlabel metal3 s 2715 353 2813 451 4 vdd
port 82 nsew
rlabel metal3 s 1392 2716 1490 2814 4 vdd
port 82 nsew
rlabel metal4 s 9902 -33 9968 25313 4 vdd
port 82 nsew
rlabel metal3 s 2715 3513 2813 3611 4 vdd
port 82 nsew
rlabel metal4 s 5926 -33 5992 25341 4 vdd
port 82 nsew
rlabel metal3 s 3094 5876 3192 5974 4 gnd
port 84 nsew
rlabel metal3 s 3094 1136 3192 1234 4 gnd
port 84 nsew
rlabel metal3 s 996 5086 1094 5184 4 gnd
port 84 nsew
rlabel metal3 s 3094 346 3192 444 4 gnd
port 84 nsew
rlabel metal4 s 5022 -33 5088 25341 4 gnd
port 84 nsew
rlabel metal4 s 7586 -63 7652 25343 4 gnd
port 84 nsew
rlabel metal3 s 2290 353 2388 451 4 gnd
port 84 nsew
rlabel metal4 s 6270 -33 6336 25341 4 gnd
port 84 nsew
rlabel metal3 s 3094 3506 3192 3604 4 gnd
port 84 nsew
rlabel metal3 s 2290 2723 2388 2821 4 gnd
port 84 nsew
rlabel metal3 s 2290 5093 2388 5191 4 gnd
port 84 nsew
rlabel metal3 s 3094 5086 3192 5184 4 gnd
port 84 nsew
rlabel metal4 s 8654 -33 8720 25313 4 gnd
port 84 nsew
rlabel metal3 s 2290 3513 2388 3611 4 gnd
port 84 nsew
rlabel metal3 s 996 2716 1094 2814 4 gnd
port 84 nsew
rlabel metal3 s 3094 2716 3192 2814 4 gnd
port 84 nsew
rlabel metal3 s 2290 5883 2388 5981 4 gnd
port 84 nsew
rlabel metal3 s 996 346 1094 444 4 gnd
port 84 nsew
rlabel metal3 s 2290 1143 2388 1241 4 gnd
port 84 nsew
<< properties >>
string FIXED_BBOX 7423 -332 7481 -331
<< end >>
