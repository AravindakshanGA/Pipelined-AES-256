magic
tech sky130A
magscale 1 2
timestamp 1543373562
<< checkpaint >>
rect -1286 -1286 22502 27356
<< metal1 >>
rect 366 25754 402 26095
rect 846 25754 882 26095
rect 1614 25754 1650 26095
rect 2094 25754 2130 26095
rect 2862 25754 2898 26095
rect 3342 25754 3378 26095
rect 4110 25754 4146 26095
rect 4590 25754 4626 26095
rect 5358 25754 5394 26095
rect 5838 25754 5874 26095
rect 6606 25754 6642 26095
rect 7086 25754 7122 26095
rect 7854 25754 7890 26095
rect 8334 25754 8370 26095
rect 9102 25754 9138 26095
rect 9582 25754 9618 26095
rect 10350 25754 10386 26095
rect 10830 25754 10866 26095
rect 11598 25754 11634 26095
rect 12078 25754 12114 26095
rect 12846 25754 12882 26095
rect 13326 25754 13362 26095
rect 14094 25754 14130 26095
rect 14574 25754 14610 26095
rect 15342 25754 15378 26095
rect 15822 25754 15858 26095
rect 16590 25754 16626 26095
rect 17070 25754 17106 26095
rect 17838 25754 17874 26095
rect 18318 25754 18354 26095
rect 19086 25754 19122 26095
rect 19566 25754 19602 26095
rect 20334 25754 20370 26095
rect 20814 25754 20850 26095
rect 366 24964 402 25596
rect 846 24964 882 25596
rect 1614 24964 1650 25596
rect 2094 24964 2130 25596
rect 2862 24964 2898 25596
rect 3342 24964 3378 25596
rect 4110 24964 4146 25596
rect 4590 24964 4626 25596
rect 5358 24964 5394 25596
rect 5838 24964 5874 25596
rect 6606 24964 6642 25596
rect 7086 24964 7122 25596
rect 7854 24964 7890 25596
rect 8334 24964 8370 25596
rect 9102 24964 9138 25596
rect 9582 24964 9618 25596
rect 10350 24964 10386 25596
rect 10830 24964 10866 25596
rect 11598 24964 11634 25596
rect 12078 24964 12114 25596
rect 12846 24964 12882 25596
rect 13326 24964 13362 25596
rect 14094 24964 14130 25596
rect 14574 24964 14610 25596
rect 15342 24964 15378 25596
rect 15822 24964 15858 25596
rect 16590 24964 16626 25596
rect 17070 24964 17106 25596
rect 17838 24964 17874 25596
rect 18318 24964 18354 25596
rect 19086 24964 19122 25596
rect 19566 24964 19602 25596
rect 20334 24964 20370 25596
rect 20814 24964 20850 25596
rect 366 24174 402 24806
rect 846 24174 882 24806
rect 1614 24174 1650 24806
rect 2094 24174 2130 24806
rect 2862 24174 2898 24806
rect 3342 24174 3378 24806
rect 4110 24174 4146 24806
rect 4590 24174 4626 24806
rect 5358 24174 5394 24806
rect 5838 24174 5874 24806
rect 6606 24174 6642 24806
rect 7086 24174 7122 24806
rect 7854 24174 7890 24806
rect 8334 24174 8370 24806
rect 9102 24174 9138 24806
rect 9582 24174 9618 24806
rect 10350 24174 10386 24806
rect 10830 24174 10866 24806
rect 11598 24174 11634 24806
rect 12078 24174 12114 24806
rect 12846 24174 12882 24806
rect 13326 24174 13362 24806
rect 14094 24174 14130 24806
rect 14574 24174 14610 24806
rect 15342 24174 15378 24806
rect 15822 24174 15858 24806
rect 16590 24174 16626 24806
rect 17070 24174 17106 24806
rect 17838 24174 17874 24806
rect 18318 24174 18354 24806
rect 19086 24174 19122 24806
rect 19566 24174 19602 24806
rect 20334 24174 20370 24806
rect 20814 24174 20850 24806
rect 366 23384 402 24016
rect 846 23384 882 24016
rect 1614 23384 1650 24016
rect 2094 23384 2130 24016
rect 2862 23384 2898 24016
rect 3342 23384 3378 24016
rect 4110 23384 4146 24016
rect 4590 23384 4626 24016
rect 5358 23384 5394 24016
rect 5838 23384 5874 24016
rect 6606 23384 6642 24016
rect 7086 23384 7122 24016
rect 7854 23384 7890 24016
rect 8334 23384 8370 24016
rect 9102 23384 9138 24016
rect 9582 23384 9618 24016
rect 10350 23384 10386 24016
rect 10830 23384 10866 24016
rect 11598 23384 11634 24016
rect 12078 23384 12114 24016
rect 12846 23384 12882 24016
rect 13326 23384 13362 24016
rect 14094 23384 14130 24016
rect 14574 23384 14610 24016
rect 15342 23384 15378 24016
rect 15822 23384 15858 24016
rect 16590 23384 16626 24016
rect 17070 23384 17106 24016
rect 17838 23384 17874 24016
rect 18318 23384 18354 24016
rect 19086 23384 19122 24016
rect 19566 23384 19602 24016
rect 20334 23384 20370 24016
rect 20814 23384 20850 24016
rect 366 22594 402 23226
rect 846 22594 882 23226
rect 1614 22594 1650 23226
rect 2094 22594 2130 23226
rect 2862 22594 2898 23226
rect 3342 22594 3378 23226
rect 4110 22594 4146 23226
rect 4590 22594 4626 23226
rect 5358 22594 5394 23226
rect 5838 22594 5874 23226
rect 6606 22594 6642 23226
rect 7086 22594 7122 23226
rect 7854 22594 7890 23226
rect 8334 22594 8370 23226
rect 9102 22594 9138 23226
rect 9582 22594 9618 23226
rect 10350 22594 10386 23226
rect 10830 22594 10866 23226
rect 11598 22594 11634 23226
rect 12078 22594 12114 23226
rect 12846 22594 12882 23226
rect 13326 22594 13362 23226
rect 14094 22594 14130 23226
rect 14574 22594 14610 23226
rect 15342 22594 15378 23226
rect 15822 22594 15858 23226
rect 16590 22594 16626 23226
rect 17070 22594 17106 23226
rect 17838 22594 17874 23226
rect 18318 22594 18354 23226
rect 19086 22594 19122 23226
rect 19566 22594 19602 23226
rect 20334 22594 20370 23226
rect 20814 22594 20850 23226
rect 366 21804 402 22436
rect 846 21804 882 22436
rect 1614 21804 1650 22436
rect 2094 21804 2130 22436
rect 2862 21804 2898 22436
rect 3342 21804 3378 22436
rect 4110 21804 4146 22436
rect 4590 21804 4626 22436
rect 5358 21804 5394 22436
rect 5838 21804 5874 22436
rect 6606 21804 6642 22436
rect 7086 21804 7122 22436
rect 7854 21804 7890 22436
rect 8334 21804 8370 22436
rect 9102 21804 9138 22436
rect 9582 21804 9618 22436
rect 10350 21804 10386 22436
rect 10830 21804 10866 22436
rect 11598 21804 11634 22436
rect 12078 21804 12114 22436
rect 12846 21804 12882 22436
rect 13326 21804 13362 22436
rect 14094 21804 14130 22436
rect 14574 21804 14610 22436
rect 15342 21804 15378 22436
rect 15822 21804 15858 22436
rect 16590 21804 16626 22436
rect 17070 21804 17106 22436
rect 17838 21804 17874 22436
rect 18318 21804 18354 22436
rect 19086 21804 19122 22436
rect 19566 21804 19602 22436
rect 20334 21804 20370 22436
rect 20814 21804 20850 22436
rect 366 21014 402 21646
rect 846 21014 882 21646
rect 1614 21014 1650 21646
rect 2094 21014 2130 21646
rect 2862 21014 2898 21646
rect 3342 21014 3378 21646
rect 4110 21014 4146 21646
rect 4590 21014 4626 21646
rect 5358 21014 5394 21646
rect 5838 21014 5874 21646
rect 6606 21014 6642 21646
rect 7086 21014 7122 21646
rect 7854 21014 7890 21646
rect 8334 21014 8370 21646
rect 9102 21014 9138 21646
rect 9582 21014 9618 21646
rect 10350 21014 10386 21646
rect 10830 21014 10866 21646
rect 11598 21014 11634 21646
rect 12078 21014 12114 21646
rect 12846 21014 12882 21646
rect 13326 21014 13362 21646
rect 14094 21014 14130 21646
rect 14574 21014 14610 21646
rect 15342 21014 15378 21646
rect 15822 21014 15858 21646
rect 16590 21014 16626 21646
rect 17070 21014 17106 21646
rect 17838 21014 17874 21646
rect 18318 21014 18354 21646
rect 19086 21014 19122 21646
rect 19566 21014 19602 21646
rect 20334 21014 20370 21646
rect 20814 21014 20850 21646
rect 366 20224 402 20856
rect 846 20224 882 20856
rect 1614 20224 1650 20856
rect 2094 20224 2130 20856
rect 2862 20224 2898 20856
rect 3342 20224 3378 20856
rect 4110 20224 4146 20856
rect 4590 20224 4626 20856
rect 5358 20224 5394 20856
rect 5838 20224 5874 20856
rect 6606 20224 6642 20856
rect 7086 20224 7122 20856
rect 7854 20224 7890 20856
rect 8334 20224 8370 20856
rect 9102 20224 9138 20856
rect 9582 20224 9618 20856
rect 10350 20224 10386 20856
rect 10830 20224 10866 20856
rect 11598 20224 11634 20856
rect 12078 20224 12114 20856
rect 12846 20224 12882 20856
rect 13326 20224 13362 20856
rect 14094 20224 14130 20856
rect 14574 20224 14610 20856
rect 15342 20224 15378 20856
rect 15822 20224 15858 20856
rect 16590 20224 16626 20856
rect 17070 20224 17106 20856
rect 17838 20224 17874 20856
rect 18318 20224 18354 20856
rect 19086 20224 19122 20856
rect 19566 20224 19602 20856
rect 20334 20224 20370 20856
rect 20814 20224 20850 20856
rect 366 19434 402 20066
rect 846 19434 882 20066
rect 1614 19434 1650 20066
rect 2094 19434 2130 20066
rect 2862 19434 2898 20066
rect 3342 19434 3378 20066
rect 4110 19434 4146 20066
rect 4590 19434 4626 20066
rect 5358 19434 5394 20066
rect 5838 19434 5874 20066
rect 6606 19434 6642 20066
rect 7086 19434 7122 20066
rect 7854 19434 7890 20066
rect 8334 19434 8370 20066
rect 9102 19434 9138 20066
rect 9582 19434 9618 20066
rect 10350 19434 10386 20066
rect 10830 19434 10866 20066
rect 11598 19434 11634 20066
rect 12078 19434 12114 20066
rect 12846 19434 12882 20066
rect 13326 19434 13362 20066
rect 14094 19434 14130 20066
rect 14574 19434 14610 20066
rect 15342 19434 15378 20066
rect 15822 19434 15858 20066
rect 16590 19434 16626 20066
rect 17070 19434 17106 20066
rect 17838 19434 17874 20066
rect 18318 19434 18354 20066
rect 19086 19434 19122 20066
rect 19566 19434 19602 20066
rect 20334 19434 20370 20066
rect 20814 19434 20850 20066
rect 366 18644 402 19276
rect 846 18644 882 19276
rect 1614 18644 1650 19276
rect 2094 18644 2130 19276
rect 2862 18644 2898 19276
rect 3342 18644 3378 19276
rect 4110 18644 4146 19276
rect 4590 18644 4626 19276
rect 5358 18644 5394 19276
rect 5838 18644 5874 19276
rect 6606 18644 6642 19276
rect 7086 18644 7122 19276
rect 7854 18644 7890 19276
rect 8334 18644 8370 19276
rect 9102 18644 9138 19276
rect 9582 18644 9618 19276
rect 10350 18644 10386 19276
rect 10830 18644 10866 19276
rect 11598 18644 11634 19276
rect 12078 18644 12114 19276
rect 12846 18644 12882 19276
rect 13326 18644 13362 19276
rect 14094 18644 14130 19276
rect 14574 18644 14610 19276
rect 15342 18644 15378 19276
rect 15822 18644 15858 19276
rect 16590 18644 16626 19276
rect 17070 18644 17106 19276
rect 17838 18644 17874 19276
rect 18318 18644 18354 19276
rect 19086 18644 19122 19276
rect 19566 18644 19602 19276
rect 20334 18644 20370 19276
rect 20814 18644 20850 19276
rect 366 17854 402 18486
rect 846 17854 882 18486
rect 1614 17854 1650 18486
rect 2094 17854 2130 18486
rect 2862 17854 2898 18486
rect 3342 17854 3378 18486
rect 4110 17854 4146 18486
rect 4590 17854 4626 18486
rect 5358 17854 5394 18486
rect 5838 17854 5874 18486
rect 6606 17854 6642 18486
rect 7086 17854 7122 18486
rect 7854 17854 7890 18486
rect 8334 17854 8370 18486
rect 9102 17854 9138 18486
rect 9582 17854 9618 18486
rect 10350 17854 10386 18486
rect 10830 17854 10866 18486
rect 11598 17854 11634 18486
rect 12078 17854 12114 18486
rect 12846 17854 12882 18486
rect 13326 17854 13362 18486
rect 14094 17854 14130 18486
rect 14574 17854 14610 18486
rect 15342 17854 15378 18486
rect 15822 17854 15858 18486
rect 16590 17854 16626 18486
rect 17070 17854 17106 18486
rect 17838 17854 17874 18486
rect 18318 17854 18354 18486
rect 19086 17854 19122 18486
rect 19566 17854 19602 18486
rect 20334 17854 20370 18486
rect 20814 17854 20850 18486
rect 366 17064 402 17696
rect 846 17064 882 17696
rect 1614 17064 1650 17696
rect 2094 17064 2130 17696
rect 2862 17064 2898 17696
rect 3342 17064 3378 17696
rect 4110 17064 4146 17696
rect 4590 17064 4626 17696
rect 5358 17064 5394 17696
rect 5838 17064 5874 17696
rect 6606 17064 6642 17696
rect 7086 17064 7122 17696
rect 7854 17064 7890 17696
rect 8334 17064 8370 17696
rect 9102 17064 9138 17696
rect 9582 17064 9618 17696
rect 10350 17064 10386 17696
rect 10830 17064 10866 17696
rect 11598 17064 11634 17696
rect 12078 17064 12114 17696
rect 12846 17064 12882 17696
rect 13326 17064 13362 17696
rect 14094 17064 14130 17696
rect 14574 17064 14610 17696
rect 15342 17064 15378 17696
rect 15822 17064 15858 17696
rect 16590 17064 16626 17696
rect 17070 17064 17106 17696
rect 17838 17064 17874 17696
rect 18318 17064 18354 17696
rect 19086 17064 19122 17696
rect 19566 17064 19602 17696
rect 20334 17064 20370 17696
rect 20814 17064 20850 17696
rect 366 16274 402 16906
rect 846 16274 882 16906
rect 1614 16274 1650 16906
rect 2094 16274 2130 16906
rect 2862 16274 2898 16906
rect 3342 16274 3378 16906
rect 4110 16274 4146 16906
rect 4590 16274 4626 16906
rect 5358 16274 5394 16906
rect 5838 16274 5874 16906
rect 6606 16274 6642 16906
rect 7086 16274 7122 16906
rect 7854 16274 7890 16906
rect 8334 16274 8370 16906
rect 9102 16274 9138 16906
rect 9582 16274 9618 16906
rect 10350 16274 10386 16906
rect 10830 16274 10866 16906
rect 11598 16274 11634 16906
rect 12078 16274 12114 16906
rect 12846 16274 12882 16906
rect 13326 16274 13362 16906
rect 14094 16274 14130 16906
rect 14574 16274 14610 16906
rect 15342 16274 15378 16906
rect 15822 16274 15858 16906
rect 16590 16274 16626 16906
rect 17070 16274 17106 16906
rect 17838 16274 17874 16906
rect 18318 16274 18354 16906
rect 19086 16274 19122 16906
rect 19566 16274 19602 16906
rect 20334 16274 20370 16906
rect 20814 16274 20850 16906
rect 366 15484 402 16116
rect 846 15484 882 16116
rect 1614 15484 1650 16116
rect 2094 15484 2130 16116
rect 2862 15484 2898 16116
rect 3342 15484 3378 16116
rect 4110 15484 4146 16116
rect 4590 15484 4626 16116
rect 5358 15484 5394 16116
rect 5838 15484 5874 16116
rect 6606 15484 6642 16116
rect 7086 15484 7122 16116
rect 7854 15484 7890 16116
rect 8334 15484 8370 16116
rect 9102 15484 9138 16116
rect 9582 15484 9618 16116
rect 10350 15484 10386 16116
rect 10830 15484 10866 16116
rect 11598 15484 11634 16116
rect 12078 15484 12114 16116
rect 12846 15484 12882 16116
rect 13326 15484 13362 16116
rect 14094 15484 14130 16116
rect 14574 15484 14610 16116
rect 15342 15484 15378 16116
rect 15822 15484 15858 16116
rect 16590 15484 16626 16116
rect 17070 15484 17106 16116
rect 17838 15484 17874 16116
rect 18318 15484 18354 16116
rect 19086 15484 19122 16116
rect 19566 15484 19602 16116
rect 20334 15484 20370 16116
rect 20814 15484 20850 16116
rect 366 14694 402 15326
rect 846 14694 882 15326
rect 1614 14694 1650 15326
rect 2094 14694 2130 15326
rect 2862 14694 2898 15326
rect 3342 14694 3378 15326
rect 4110 14694 4146 15326
rect 4590 14694 4626 15326
rect 5358 14694 5394 15326
rect 5838 14694 5874 15326
rect 6606 14694 6642 15326
rect 7086 14694 7122 15326
rect 7854 14694 7890 15326
rect 8334 14694 8370 15326
rect 9102 14694 9138 15326
rect 9582 14694 9618 15326
rect 10350 14694 10386 15326
rect 10830 14694 10866 15326
rect 11598 14694 11634 15326
rect 12078 14694 12114 15326
rect 12846 14694 12882 15326
rect 13326 14694 13362 15326
rect 14094 14694 14130 15326
rect 14574 14694 14610 15326
rect 15342 14694 15378 15326
rect 15822 14694 15858 15326
rect 16590 14694 16626 15326
rect 17070 14694 17106 15326
rect 17838 14694 17874 15326
rect 18318 14694 18354 15326
rect 19086 14694 19122 15326
rect 19566 14694 19602 15326
rect 20334 14694 20370 15326
rect 20814 14694 20850 15326
rect 366 13904 402 14536
rect 846 13904 882 14536
rect 1614 13904 1650 14536
rect 2094 13904 2130 14536
rect 2862 13904 2898 14536
rect 3342 13904 3378 14536
rect 4110 13904 4146 14536
rect 4590 13904 4626 14536
rect 5358 13904 5394 14536
rect 5838 13904 5874 14536
rect 6606 13904 6642 14536
rect 7086 13904 7122 14536
rect 7854 13904 7890 14536
rect 8334 13904 8370 14536
rect 9102 13904 9138 14536
rect 9582 13904 9618 14536
rect 10350 13904 10386 14536
rect 10830 13904 10866 14536
rect 11598 13904 11634 14536
rect 12078 13904 12114 14536
rect 12846 13904 12882 14536
rect 13326 13904 13362 14536
rect 14094 13904 14130 14536
rect 14574 13904 14610 14536
rect 15342 13904 15378 14536
rect 15822 13904 15858 14536
rect 16590 13904 16626 14536
rect 17070 13904 17106 14536
rect 17838 13904 17874 14536
rect 18318 13904 18354 14536
rect 19086 13904 19122 14536
rect 19566 13904 19602 14536
rect 20334 13904 20370 14536
rect 20814 13904 20850 14536
rect 366 13114 402 13746
rect 846 13114 882 13746
rect 1614 13114 1650 13746
rect 2094 13114 2130 13746
rect 2862 13114 2898 13746
rect 3342 13114 3378 13746
rect 4110 13114 4146 13746
rect 4590 13114 4626 13746
rect 5358 13114 5394 13746
rect 5838 13114 5874 13746
rect 6606 13114 6642 13746
rect 7086 13114 7122 13746
rect 7854 13114 7890 13746
rect 8334 13114 8370 13746
rect 9102 13114 9138 13746
rect 9582 13114 9618 13746
rect 10350 13114 10386 13746
rect 10830 13114 10866 13746
rect 11598 13114 11634 13746
rect 12078 13114 12114 13746
rect 12846 13114 12882 13746
rect 13326 13114 13362 13746
rect 14094 13114 14130 13746
rect 14574 13114 14610 13746
rect 15342 13114 15378 13746
rect 15822 13114 15858 13746
rect 16590 13114 16626 13746
rect 17070 13114 17106 13746
rect 17838 13114 17874 13746
rect 18318 13114 18354 13746
rect 19086 13114 19122 13746
rect 19566 13114 19602 13746
rect 20334 13114 20370 13746
rect 20814 13114 20850 13746
rect 366 12324 402 12956
rect 846 12324 882 12956
rect 1614 12324 1650 12956
rect 2094 12324 2130 12956
rect 2862 12324 2898 12956
rect 3342 12324 3378 12956
rect 4110 12324 4146 12956
rect 4590 12324 4626 12956
rect 5358 12324 5394 12956
rect 5838 12324 5874 12956
rect 6606 12324 6642 12956
rect 7086 12324 7122 12956
rect 7854 12324 7890 12956
rect 8334 12324 8370 12956
rect 9102 12324 9138 12956
rect 9582 12324 9618 12956
rect 10350 12324 10386 12956
rect 10830 12324 10866 12956
rect 11598 12324 11634 12956
rect 12078 12324 12114 12956
rect 12846 12324 12882 12956
rect 13326 12324 13362 12956
rect 14094 12324 14130 12956
rect 14574 12324 14610 12956
rect 15342 12324 15378 12956
rect 15822 12324 15858 12956
rect 16590 12324 16626 12956
rect 17070 12324 17106 12956
rect 17838 12324 17874 12956
rect 18318 12324 18354 12956
rect 19086 12324 19122 12956
rect 19566 12324 19602 12956
rect 20334 12324 20370 12956
rect 20814 12324 20850 12956
rect 366 11534 402 12166
rect 846 11534 882 12166
rect 1614 11534 1650 12166
rect 2094 11534 2130 12166
rect 2862 11534 2898 12166
rect 3342 11534 3378 12166
rect 4110 11534 4146 12166
rect 4590 11534 4626 12166
rect 5358 11534 5394 12166
rect 5838 11534 5874 12166
rect 6606 11534 6642 12166
rect 7086 11534 7122 12166
rect 7854 11534 7890 12166
rect 8334 11534 8370 12166
rect 9102 11534 9138 12166
rect 9582 11534 9618 12166
rect 10350 11534 10386 12166
rect 10830 11534 10866 12166
rect 11598 11534 11634 12166
rect 12078 11534 12114 12166
rect 12846 11534 12882 12166
rect 13326 11534 13362 12166
rect 14094 11534 14130 12166
rect 14574 11534 14610 12166
rect 15342 11534 15378 12166
rect 15822 11534 15858 12166
rect 16590 11534 16626 12166
rect 17070 11534 17106 12166
rect 17838 11534 17874 12166
rect 18318 11534 18354 12166
rect 19086 11534 19122 12166
rect 19566 11534 19602 12166
rect 20334 11534 20370 12166
rect 20814 11534 20850 12166
rect 366 10744 402 11376
rect 846 10744 882 11376
rect 1614 10744 1650 11376
rect 2094 10744 2130 11376
rect 2862 10744 2898 11376
rect 3342 10744 3378 11376
rect 4110 10744 4146 11376
rect 4590 10744 4626 11376
rect 5358 10744 5394 11376
rect 5838 10744 5874 11376
rect 6606 10744 6642 11376
rect 7086 10744 7122 11376
rect 7854 10744 7890 11376
rect 8334 10744 8370 11376
rect 9102 10744 9138 11376
rect 9582 10744 9618 11376
rect 10350 10744 10386 11376
rect 10830 10744 10866 11376
rect 11598 10744 11634 11376
rect 12078 10744 12114 11376
rect 12846 10744 12882 11376
rect 13326 10744 13362 11376
rect 14094 10744 14130 11376
rect 14574 10744 14610 11376
rect 15342 10744 15378 11376
rect 15822 10744 15858 11376
rect 16590 10744 16626 11376
rect 17070 10744 17106 11376
rect 17838 10744 17874 11376
rect 18318 10744 18354 11376
rect 19086 10744 19122 11376
rect 19566 10744 19602 11376
rect 20334 10744 20370 11376
rect 20814 10744 20850 11376
rect 366 9954 402 10586
rect 846 9954 882 10586
rect 1614 9954 1650 10586
rect 2094 9954 2130 10586
rect 2862 9954 2898 10586
rect 3342 9954 3378 10586
rect 4110 9954 4146 10586
rect 4590 9954 4626 10586
rect 5358 9954 5394 10586
rect 5838 9954 5874 10586
rect 6606 9954 6642 10586
rect 7086 9954 7122 10586
rect 7854 9954 7890 10586
rect 8334 9954 8370 10586
rect 9102 9954 9138 10586
rect 9582 9954 9618 10586
rect 10350 9954 10386 10586
rect 10830 9954 10866 10586
rect 11598 9954 11634 10586
rect 12078 9954 12114 10586
rect 12846 9954 12882 10586
rect 13326 9954 13362 10586
rect 14094 9954 14130 10586
rect 14574 9954 14610 10586
rect 15342 9954 15378 10586
rect 15822 9954 15858 10586
rect 16590 9954 16626 10586
rect 17070 9954 17106 10586
rect 17838 9954 17874 10586
rect 18318 9954 18354 10586
rect 19086 9954 19122 10586
rect 19566 9954 19602 10586
rect 20334 9954 20370 10586
rect 20814 9954 20850 10586
rect 366 9164 402 9796
rect 846 9164 882 9796
rect 1614 9164 1650 9796
rect 2094 9164 2130 9796
rect 2862 9164 2898 9796
rect 3342 9164 3378 9796
rect 4110 9164 4146 9796
rect 4590 9164 4626 9796
rect 5358 9164 5394 9796
rect 5838 9164 5874 9796
rect 6606 9164 6642 9796
rect 7086 9164 7122 9796
rect 7854 9164 7890 9796
rect 8334 9164 8370 9796
rect 9102 9164 9138 9796
rect 9582 9164 9618 9796
rect 10350 9164 10386 9796
rect 10830 9164 10866 9796
rect 11598 9164 11634 9796
rect 12078 9164 12114 9796
rect 12846 9164 12882 9796
rect 13326 9164 13362 9796
rect 14094 9164 14130 9796
rect 14574 9164 14610 9796
rect 15342 9164 15378 9796
rect 15822 9164 15858 9796
rect 16590 9164 16626 9796
rect 17070 9164 17106 9796
rect 17838 9164 17874 9796
rect 18318 9164 18354 9796
rect 19086 9164 19122 9796
rect 19566 9164 19602 9796
rect 20334 9164 20370 9796
rect 20814 9164 20850 9796
rect 366 8374 402 9006
rect 846 8374 882 9006
rect 1614 8374 1650 9006
rect 2094 8374 2130 9006
rect 2862 8374 2898 9006
rect 3342 8374 3378 9006
rect 4110 8374 4146 9006
rect 4590 8374 4626 9006
rect 5358 8374 5394 9006
rect 5838 8374 5874 9006
rect 6606 8374 6642 9006
rect 7086 8374 7122 9006
rect 7854 8374 7890 9006
rect 8334 8374 8370 9006
rect 9102 8374 9138 9006
rect 9582 8374 9618 9006
rect 10350 8374 10386 9006
rect 10830 8374 10866 9006
rect 11598 8374 11634 9006
rect 12078 8374 12114 9006
rect 12846 8374 12882 9006
rect 13326 8374 13362 9006
rect 14094 8374 14130 9006
rect 14574 8374 14610 9006
rect 15342 8374 15378 9006
rect 15822 8374 15858 9006
rect 16590 8374 16626 9006
rect 17070 8374 17106 9006
rect 17838 8374 17874 9006
rect 18318 8374 18354 9006
rect 19086 8374 19122 9006
rect 19566 8374 19602 9006
rect 20334 8374 20370 9006
rect 20814 8374 20850 9006
rect 366 7584 402 8216
rect 846 7584 882 8216
rect 1614 7584 1650 8216
rect 2094 7584 2130 8216
rect 2862 7584 2898 8216
rect 3342 7584 3378 8216
rect 4110 7584 4146 8216
rect 4590 7584 4626 8216
rect 5358 7584 5394 8216
rect 5838 7584 5874 8216
rect 6606 7584 6642 8216
rect 7086 7584 7122 8216
rect 7854 7584 7890 8216
rect 8334 7584 8370 8216
rect 9102 7584 9138 8216
rect 9582 7584 9618 8216
rect 10350 7584 10386 8216
rect 10830 7584 10866 8216
rect 11598 7584 11634 8216
rect 12078 7584 12114 8216
rect 12846 7584 12882 8216
rect 13326 7584 13362 8216
rect 14094 7584 14130 8216
rect 14574 7584 14610 8216
rect 15342 7584 15378 8216
rect 15822 7584 15858 8216
rect 16590 7584 16626 8216
rect 17070 7584 17106 8216
rect 17838 7584 17874 8216
rect 18318 7584 18354 8216
rect 19086 7584 19122 8216
rect 19566 7584 19602 8216
rect 20334 7584 20370 8216
rect 20814 7584 20850 8216
rect 366 6794 402 7426
rect 846 6794 882 7426
rect 1614 6794 1650 7426
rect 2094 6794 2130 7426
rect 2862 6794 2898 7426
rect 3342 6794 3378 7426
rect 4110 6794 4146 7426
rect 4590 6794 4626 7426
rect 5358 6794 5394 7426
rect 5838 6794 5874 7426
rect 6606 6794 6642 7426
rect 7086 6794 7122 7426
rect 7854 6794 7890 7426
rect 8334 6794 8370 7426
rect 9102 6794 9138 7426
rect 9582 6794 9618 7426
rect 10350 6794 10386 7426
rect 10830 6794 10866 7426
rect 11598 6794 11634 7426
rect 12078 6794 12114 7426
rect 12846 6794 12882 7426
rect 13326 6794 13362 7426
rect 14094 6794 14130 7426
rect 14574 6794 14610 7426
rect 15342 6794 15378 7426
rect 15822 6794 15858 7426
rect 16590 6794 16626 7426
rect 17070 6794 17106 7426
rect 17838 6794 17874 7426
rect 18318 6794 18354 7426
rect 19086 6794 19122 7426
rect 19566 6794 19602 7426
rect 20334 6794 20370 7426
rect 20814 6794 20850 7426
rect 366 6004 402 6636
rect 846 6004 882 6636
rect 1614 6004 1650 6636
rect 2094 6004 2130 6636
rect 2862 6004 2898 6636
rect 3342 6004 3378 6636
rect 4110 6004 4146 6636
rect 4590 6004 4626 6636
rect 5358 6004 5394 6636
rect 5838 6004 5874 6636
rect 6606 6004 6642 6636
rect 7086 6004 7122 6636
rect 7854 6004 7890 6636
rect 8334 6004 8370 6636
rect 9102 6004 9138 6636
rect 9582 6004 9618 6636
rect 10350 6004 10386 6636
rect 10830 6004 10866 6636
rect 11598 6004 11634 6636
rect 12078 6004 12114 6636
rect 12846 6004 12882 6636
rect 13326 6004 13362 6636
rect 14094 6004 14130 6636
rect 14574 6004 14610 6636
rect 15342 6004 15378 6636
rect 15822 6004 15858 6636
rect 16590 6004 16626 6636
rect 17070 6004 17106 6636
rect 17838 6004 17874 6636
rect 18318 6004 18354 6636
rect 19086 6004 19122 6636
rect 19566 6004 19602 6636
rect 20334 6004 20370 6636
rect 20814 6004 20850 6636
rect 366 5214 402 5846
rect 846 5214 882 5846
rect 1614 5214 1650 5846
rect 2094 5214 2130 5846
rect 2862 5214 2898 5846
rect 3342 5214 3378 5846
rect 4110 5214 4146 5846
rect 4590 5214 4626 5846
rect 5358 5214 5394 5846
rect 5838 5214 5874 5846
rect 6606 5214 6642 5846
rect 7086 5214 7122 5846
rect 7854 5214 7890 5846
rect 8334 5214 8370 5846
rect 9102 5214 9138 5846
rect 9582 5214 9618 5846
rect 10350 5214 10386 5846
rect 10830 5214 10866 5846
rect 11598 5214 11634 5846
rect 12078 5214 12114 5846
rect 12846 5214 12882 5846
rect 13326 5214 13362 5846
rect 14094 5214 14130 5846
rect 14574 5214 14610 5846
rect 15342 5214 15378 5846
rect 15822 5214 15858 5846
rect 16590 5214 16626 5846
rect 17070 5214 17106 5846
rect 17838 5214 17874 5846
rect 18318 5214 18354 5846
rect 19086 5214 19122 5846
rect 19566 5214 19602 5846
rect 20334 5214 20370 5846
rect 20814 5214 20850 5846
rect 366 4424 402 5056
rect 846 4424 882 5056
rect 1614 4424 1650 5056
rect 2094 4424 2130 5056
rect 2862 4424 2898 5056
rect 3342 4424 3378 5056
rect 4110 4424 4146 5056
rect 4590 4424 4626 5056
rect 5358 4424 5394 5056
rect 5838 4424 5874 5056
rect 6606 4424 6642 5056
rect 7086 4424 7122 5056
rect 7854 4424 7890 5056
rect 8334 4424 8370 5056
rect 9102 4424 9138 5056
rect 9582 4424 9618 5056
rect 10350 4424 10386 5056
rect 10830 4424 10866 5056
rect 11598 4424 11634 5056
rect 12078 4424 12114 5056
rect 12846 4424 12882 5056
rect 13326 4424 13362 5056
rect 14094 4424 14130 5056
rect 14574 4424 14610 5056
rect 15342 4424 15378 5056
rect 15822 4424 15858 5056
rect 16590 4424 16626 5056
rect 17070 4424 17106 5056
rect 17838 4424 17874 5056
rect 18318 4424 18354 5056
rect 19086 4424 19122 5056
rect 19566 4424 19602 5056
rect 20334 4424 20370 5056
rect 20814 4424 20850 5056
rect 366 3634 402 4266
rect 846 3634 882 4266
rect 1614 3634 1650 4266
rect 2094 3634 2130 4266
rect 2862 3634 2898 4266
rect 3342 3634 3378 4266
rect 4110 3634 4146 4266
rect 4590 3634 4626 4266
rect 5358 3634 5394 4266
rect 5838 3634 5874 4266
rect 6606 3634 6642 4266
rect 7086 3634 7122 4266
rect 7854 3634 7890 4266
rect 8334 3634 8370 4266
rect 9102 3634 9138 4266
rect 9582 3634 9618 4266
rect 10350 3634 10386 4266
rect 10830 3634 10866 4266
rect 11598 3634 11634 4266
rect 12078 3634 12114 4266
rect 12846 3634 12882 4266
rect 13326 3634 13362 4266
rect 14094 3634 14130 4266
rect 14574 3634 14610 4266
rect 15342 3634 15378 4266
rect 15822 3634 15858 4266
rect 16590 3634 16626 4266
rect 17070 3634 17106 4266
rect 17838 3634 17874 4266
rect 18318 3634 18354 4266
rect 19086 3634 19122 4266
rect 19566 3634 19602 4266
rect 20334 3634 20370 4266
rect 20814 3634 20850 4266
rect 366 2844 402 3476
rect 846 2844 882 3476
rect 1614 2844 1650 3476
rect 2094 2844 2130 3476
rect 2862 2844 2898 3476
rect 3342 2844 3378 3476
rect 4110 2844 4146 3476
rect 4590 2844 4626 3476
rect 5358 2844 5394 3476
rect 5838 2844 5874 3476
rect 6606 2844 6642 3476
rect 7086 2844 7122 3476
rect 7854 2844 7890 3476
rect 8334 2844 8370 3476
rect 9102 2844 9138 3476
rect 9582 2844 9618 3476
rect 10350 2844 10386 3476
rect 10830 2844 10866 3476
rect 11598 2844 11634 3476
rect 12078 2844 12114 3476
rect 12846 2844 12882 3476
rect 13326 2844 13362 3476
rect 14094 2844 14130 3476
rect 14574 2844 14610 3476
rect 15342 2844 15378 3476
rect 15822 2844 15858 3476
rect 16590 2844 16626 3476
rect 17070 2844 17106 3476
rect 17838 2844 17874 3476
rect 18318 2844 18354 3476
rect 19086 2844 19122 3476
rect 19566 2844 19602 3476
rect 20334 2844 20370 3476
rect 20814 2844 20850 3476
rect 366 2054 402 2686
rect 846 2054 882 2686
rect 1614 2054 1650 2686
rect 2094 2054 2130 2686
rect 2862 2054 2898 2686
rect 3342 2054 3378 2686
rect 4110 2054 4146 2686
rect 4590 2054 4626 2686
rect 5358 2054 5394 2686
rect 5838 2054 5874 2686
rect 6606 2054 6642 2686
rect 7086 2054 7122 2686
rect 7854 2054 7890 2686
rect 8334 2054 8370 2686
rect 9102 2054 9138 2686
rect 9582 2054 9618 2686
rect 10350 2054 10386 2686
rect 10830 2054 10866 2686
rect 11598 2054 11634 2686
rect 12078 2054 12114 2686
rect 12846 2054 12882 2686
rect 13326 2054 13362 2686
rect 14094 2054 14130 2686
rect 14574 2054 14610 2686
rect 15342 2054 15378 2686
rect 15822 2054 15858 2686
rect 16590 2054 16626 2686
rect 17070 2054 17106 2686
rect 17838 2054 17874 2686
rect 18318 2054 18354 2686
rect 19086 2054 19122 2686
rect 19566 2054 19602 2686
rect 20334 2054 20370 2686
rect 20814 2054 20850 2686
rect 366 1264 402 1896
rect 846 1264 882 1896
rect 1614 1264 1650 1896
rect 2094 1264 2130 1896
rect 2862 1264 2898 1896
rect 3342 1264 3378 1896
rect 4110 1264 4146 1896
rect 4590 1264 4626 1896
rect 5358 1264 5394 1896
rect 5838 1264 5874 1896
rect 6606 1264 6642 1896
rect 7086 1264 7122 1896
rect 7854 1264 7890 1896
rect 8334 1264 8370 1896
rect 9102 1264 9138 1896
rect 9582 1264 9618 1896
rect 10350 1264 10386 1896
rect 10830 1264 10866 1896
rect 11598 1264 11634 1896
rect 12078 1264 12114 1896
rect 12846 1264 12882 1896
rect 13326 1264 13362 1896
rect 14094 1264 14130 1896
rect 14574 1264 14610 1896
rect 15342 1264 15378 1896
rect 15822 1264 15858 1896
rect 16590 1264 16626 1896
rect 17070 1264 17106 1896
rect 17838 1264 17874 1896
rect 18318 1264 18354 1896
rect 19086 1264 19122 1896
rect 19566 1264 19602 1896
rect 20334 1264 20370 1896
rect 20814 1264 20850 1896
rect 366 474 402 1106
rect 846 474 882 1106
rect 1614 474 1650 1106
rect 2094 474 2130 1106
rect 2862 474 2898 1106
rect 3342 474 3378 1106
rect 4110 474 4146 1106
rect 4590 474 4626 1106
rect 5358 474 5394 1106
rect 5838 474 5874 1106
rect 6606 474 6642 1106
rect 7086 474 7122 1106
rect 7854 474 7890 1106
rect 8334 474 8370 1106
rect 9102 474 9138 1106
rect 9582 474 9618 1106
rect 10350 474 10386 1106
rect 10830 474 10866 1106
rect 11598 474 11634 1106
rect 12078 474 12114 1106
rect 12846 474 12882 1106
rect 13326 474 13362 1106
rect 14094 474 14130 1106
rect 14574 474 14610 1106
rect 15342 474 15378 1106
rect 15822 474 15858 1106
rect 16590 474 16626 1106
rect 17070 474 17106 1106
rect 17838 474 17874 1106
rect 18318 474 18354 1106
rect 19086 474 19122 1106
rect 19566 474 19602 1106
rect 20334 474 20370 1106
rect 20814 474 20850 1106
rect 222 0 258 28
rect 294 0 330 28
rect 366 -25 402 316
rect 438 0 474 28
rect 510 0 546 28
rect 702 0 738 28
rect 774 0 810 28
rect 846 -25 882 316
rect 918 0 954 28
rect 990 0 1026 28
rect 1470 0 1506 28
rect 1542 0 1578 28
rect 1614 -25 1650 316
rect 1686 0 1722 28
rect 1758 0 1794 28
rect 1950 0 1986 28
rect 2022 0 2058 28
rect 2094 -25 2130 316
rect 2166 0 2202 28
rect 2238 0 2274 28
rect 2718 0 2754 28
rect 2790 0 2826 28
rect 2862 -25 2898 316
rect 2934 0 2970 28
rect 3006 0 3042 28
rect 3198 0 3234 28
rect 3270 0 3306 28
rect 3342 -25 3378 316
rect 3414 0 3450 28
rect 3486 0 3522 28
rect 3966 0 4002 28
rect 4038 0 4074 28
rect 4110 -25 4146 316
rect 4182 0 4218 28
rect 4254 0 4290 28
rect 4446 0 4482 28
rect 4518 0 4554 28
rect 4590 -25 4626 316
rect 4662 0 4698 28
rect 4734 0 4770 28
rect 5214 0 5250 28
rect 5286 0 5322 28
rect 5358 -25 5394 316
rect 5430 0 5466 28
rect 5502 0 5538 28
rect 5694 0 5730 28
rect 5766 0 5802 28
rect 5838 -25 5874 316
rect 5910 0 5946 28
rect 5982 0 6018 28
rect 6462 0 6498 28
rect 6534 0 6570 28
rect 6606 -25 6642 316
rect 6678 0 6714 28
rect 6750 0 6786 28
rect 6942 0 6978 28
rect 7014 0 7050 28
rect 7086 -25 7122 316
rect 7158 0 7194 28
rect 7230 0 7266 28
rect 7710 0 7746 28
rect 7782 0 7818 28
rect 7854 -25 7890 316
rect 7926 0 7962 28
rect 7998 0 8034 28
rect 8190 0 8226 28
rect 8262 0 8298 28
rect 8334 -25 8370 316
rect 8406 0 8442 28
rect 8478 0 8514 28
rect 8958 0 8994 28
rect 9030 0 9066 28
rect 9102 -25 9138 316
rect 9174 0 9210 28
rect 9246 0 9282 28
rect 9438 0 9474 28
rect 9510 0 9546 28
rect 9582 -25 9618 316
rect 9654 0 9690 28
rect 9726 0 9762 28
rect 10206 0 10242 28
rect 10278 0 10314 28
rect 10350 -25 10386 316
rect 10422 0 10458 28
rect 10494 0 10530 28
rect 10686 0 10722 28
rect 10758 0 10794 28
rect 10830 -25 10866 316
rect 10902 0 10938 28
rect 10974 0 11010 28
rect 11454 0 11490 28
rect 11526 0 11562 28
rect 11598 -25 11634 316
rect 11670 0 11706 28
rect 11742 0 11778 28
rect 11934 0 11970 28
rect 12006 0 12042 28
rect 12078 -25 12114 316
rect 12150 0 12186 28
rect 12222 0 12258 28
rect 12702 0 12738 28
rect 12774 0 12810 28
rect 12846 -25 12882 316
rect 12918 0 12954 28
rect 12990 0 13026 28
rect 13182 0 13218 28
rect 13254 0 13290 28
rect 13326 -25 13362 316
rect 13398 0 13434 28
rect 13470 0 13506 28
rect 13950 0 13986 28
rect 14022 0 14058 28
rect 14094 -25 14130 316
rect 14166 0 14202 28
rect 14238 0 14274 28
rect 14430 0 14466 28
rect 14502 0 14538 28
rect 14574 -25 14610 316
rect 14646 0 14682 28
rect 14718 0 14754 28
rect 15198 0 15234 28
rect 15270 0 15306 28
rect 15342 -25 15378 316
rect 15414 0 15450 28
rect 15486 0 15522 28
rect 15678 0 15714 28
rect 15750 0 15786 28
rect 15822 -25 15858 316
rect 15894 0 15930 28
rect 15966 0 16002 28
rect 16446 0 16482 28
rect 16518 0 16554 28
rect 16590 -25 16626 316
rect 16662 0 16698 28
rect 16734 0 16770 28
rect 16926 0 16962 28
rect 16998 0 17034 28
rect 17070 -25 17106 316
rect 17142 0 17178 28
rect 17214 0 17250 28
rect 17694 0 17730 28
rect 17766 0 17802 28
rect 17838 -25 17874 316
rect 17910 0 17946 28
rect 17982 0 18018 28
rect 18174 0 18210 28
rect 18246 0 18282 28
rect 18318 -25 18354 316
rect 18390 0 18426 28
rect 18462 0 18498 28
rect 18942 0 18978 28
rect 19014 0 19050 28
rect 19086 -25 19122 316
rect 19158 0 19194 28
rect 19230 0 19266 28
rect 19422 0 19458 28
rect 19494 0 19530 28
rect 19566 -25 19602 316
rect 19638 0 19674 28
rect 19710 0 19746 28
rect 20190 0 20226 28
rect 20262 0 20298 28
rect 20334 -25 20370 316
rect 20406 0 20442 28
rect 20478 0 20514 28
rect 20670 0 20706 28
rect 20742 0 20778 28
rect 20814 -25 20850 316
rect 20886 0 20922 28
rect 20958 0 20994 28
<< metal2 >>
rect 0 25998 28 26046
rect 330 25874 438 25950
rect 810 25874 918 25950
rect 1578 25874 1686 25950
rect 2058 25874 2166 25950
rect 2826 25874 2934 25950
rect 3306 25874 3414 25950
rect 4074 25874 4182 25950
rect 4554 25874 4662 25950
rect 5322 25874 5430 25950
rect 5802 25874 5910 25950
rect 6570 25874 6678 25950
rect 7050 25874 7158 25950
rect 7818 25874 7926 25950
rect 8298 25874 8406 25950
rect 9066 25874 9174 25950
rect 9546 25874 9654 25950
rect 10314 25874 10422 25950
rect 10794 25874 10902 25950
rect 11562 25874 11670 25950
rect 12042 25874 12150 25950
rect 12810 25874 12918 25950
rect 13290 25874 13398 25950
rect 14058 25874 14166 25950
rect 14538 25874 14646 25950
rect 15306 25874 15414 25950
rect 15786 25874 15894 25950
rect 16554 25874 16662 25950
rect 17034 25874 17142 25950
rect 17802 25874 17910 25950
rect 18282 25874 18390 25950
rect 19050 25874 19158 25950
rect 19530 25874 19638 25950
rect 20298 25874 20406 25950
rect 20778 25874 20886 25950
rect 0 25778 28 25826
rect 330 25620 438 25730
rect 810 25620 918 25730
rect 1578 25620 1686 25730
rect 2058 25620 2166 25730
rect 2826 25620 2934 25730
rect 3306 25620 3414 25730
rect 4074 25620 4182 25730
rect 4554 25620 4662 25730
rect 5322 25620 5430 25730
rect 5802 25620 5910 25730
rect 6570 25620 6678 25730
rect 7050 25620 7158 25730
rect 7818 25620 7926 25730
rect 8298 25620 8406 25730
rect 9066 25620 9174 25730
rect 9546 25620 9654 25730
rect 10314 25620 10422 25730
rect 10794 25620 10902 25730
rect 11562 25620 11670 25730
rect 12042 25620 12150 25730
rect 12810 25620 12918 25730
rect 13290 25620 13398 25730
rect 14058 25620 14166 25730
rect 14538 25620 14646 25730
rect 15306 25620 15414 25730
rect 15786 25620 15894 25730
rect 16554 25620 16662 25730
rect 17034 25620 17142 25730
rect 17802 25620 17910 25730
rect 18282 25620 18390 25730
rect 19050 25620 19158 25730
rect 19530 25620 19638 25730
rect 20298 25620 20406 25730
rect 20778 25620 20886 25730
rect 0 25524 28 25572
rect 330 25400 438 25476
rect 810 25400 918 25476
rect 1578 25400 1686 25476
rect 2058 25400 2166 25476
rect 2826 25400 2934 25476
rect 3306 25400 3414 25476
rect 4074 25400 4182 25476
rect 4554 25400 4662 25476
rect 5322 25400 5430 25476
rect 5802 25400 5910 25476
rect 6570 25400 6678 25476
rect 7050 25400 7158 25476
rect 7818 25400 7926 25476
rect 8298 25400 8406 25476
rect 9066 25400 9174 25476
rect 9546 25400 9654 25476
rect 10314 25400 10422 25476
rect 10794 25400 10902 25476
rect 11562 25400 11670 25476
rect 12042 25400 12150 25476
rect 12810 25400 12918 25476
rect 13290 25400 13398 25476
rect 14058 25400 14166 25476
rect 14538 25400 14646 25476
rect 15306 25400 15414 25476
rect 15786 25400 15894 25476
rect 16554 25400 16662 25476
rect 17034 25400 17142 25476
rect 17802 25400 17910 25476
rect 18282 25400 18390 25476
rect 19050 25400 19158 25476
rect 19530 25400 19638 25476
rect 20298 25400 20406 25476
rect 20778 25400 20886 25476
rect 0 25304 28 25352
rect 0 25208 28 25256
rect 330 25084 438 25160
rect 810 25084 918 25160
rect 1578 25084 1686 25160
rect 2058 25084 2166 25160
rect 2826 25084 2934 25160
rect 3306 25084 3414 25160
rect 4074 25084 4182 25160
rect 4554 25084 4662 25160
rect 5322 25084 5430 25160
rect 5802 25084 5910 25160
rect 6570 25084 6678 25160
rect 7050 25084 7158 25160
rect 7818 25084 7926 25160
rect 8298 25084 8406 25160
rect 9066 25084 9174 25160
rect 9546 25084 9654 25160
rect 10314 25084 10422 25160
rect 10794 25084 10902 25160
rect 11562 25084 11670 25160
rect 12042 25084 12150 25160
rect 12810 25084 12918 25160
rect 13290 25084 13398 25160
rect 14058 25084 14166 25160
rect 14538 25084 14646 25160
rect 15306 25084 15414 25160
rect 15786 25084 15894 25160
rect 16554 25084 16662 25160
rect 17034 25084 17142 25160
rect 17802 25084 17910 25160
rect 18282 25084 18390 25160
rect 19050 25084 19158 25160
rect 19530 25084 19638 25160
rect 20298 25084 20406 25160
rect 20778 25084 20886 25160
rect 0 24988 28 25036
rect 330 24830 438 24940
rect 810 24830 918 24940
rect 1578 24830 1686 24940
rect 2058 24830 2166 24940
rect 2826 24830 2934 24940
rect 3306 24830 3414 24940
rect 4074 24830 4182 24940
rect 4554 24830 4662 24940
rect 5322 24830 5430 24940
rect 5802 24830 5910 24940
rect 6570 24830 6678 24940
rect 7050 24830 7158 24940
rect 7818 24830 7926 24940
rect 8298 24830 8406 24940
rect 9066 24830 9174 24940
rect 9546 24830 9654 24940
rect 10314 24830 10422 24940
rect 10794 24830 10902 24940
rect 11562 24830 11670 24940
rect 12042 24830 12150 24940
rect 12810 24830 12918 24940
rect 13290 24830 13398 24940
rect 14058 24830 14166 24940
rect 14538 24830 14646 24940
rect 15306 24830 15414 24940
rect 15786 24830 15894 24940
rect 16554 24830 16662 24940
rect 17034 24830 17142 24940
rect 17802 24830 17910 24940
rect 18282 24830 18390 24940
rect 19050 24830 19158 24940
rect 19530 24830 19638 24940
rect 20298 24830 20406 24940
rect 20778 24830 20886 24940
rect 0 24734 28 24782
rect 330 24610 438 24686
rect 810 24610 918 24686
rect 1578 24610 1686 24686
rect 2058 24610 2166 24686
rect 2826 24610 2934 24686
rect 3306 24610 3414 24686
rect 4074 24610 4182 24686
rect 4554 24610 4662 24686
rect 5322 24610 5430 24686
rect 5802 24610 5910 24686
rect 6570 24610 6678 24686
rect 7050 24610 7158 24686
rect 7818 24610 7926 24686
rect 8298 24610 8406 24686
rect 9066 24610 9174 24686
rect 9546 24610 9654 24686
rect 10314 24610 10422 24686
rect 10794 24610 10902 24686
rect 11562 24610 11670 24686
rect 12042 24610 12150 24686
rect 12810 24610 12918 24686
rect 13290 24610 13398 24686
rect 14058 24610 14166 24686
rect 14538 24610 14646 24686
rect 15306 24610 15414 24686
rect 15786 24610 15894 24686
rect 16554 24610 16662 24686
rect 17034 24610 17142 24686
rect 17802 24610 17910 24686
rect 18282 24610 18390 24686
rect 19050 24610 19158 24686
rect 19530 24610 19638 24686
rect 20298 24610 20406 24686
rect 20778 24610 20886 24686
rect 0 24514 28 24562
rect 0 24418 28 24466
rect 330 24294 438 24370
rect 810 24294 918 24370
rect 1578 24294 1686 24370
rect 2058 24294 2166 24370
rect 2826 24294 2934 24370
rect 3306 24294 3414 24370
rect 4074 24294 4182 24370
rect 4554 24294 4662 24370
rect 5322 24294 5430 24370
rect 5802 24294 5910 24370
rect 6570 24294 6678 24370
rect 7050 24294 7158 24370
rect 7818 24294 7926 24370
rect 8298 24294 8406 24370
rect 9066 24294 9174 24370
rect 9546 24294 9654 24370
rect 10314 24294 10422 24370
rect 10794 24294 10902 24370
rect 11562 24294 11670 24370
rect 12042 24294 12150 24370
rect 12810 24294 12918 24370
rect 13290 24294 13398 24370
rect 14058 24294 14166 24370
rect 14538 24294 14646 24370
rect 15306 24294 15414 24370
rect 15786 24294 15894 24370
rect 16554 24294 16662 24370
rect 17034 24294 17142 24370
rect 17802 24294 17910 24370
rect 18282 24294 18390 24370
rect 19050 24294 19158 24370
rect 19530 24294 19638 24370
rect 20298 24294 20406 24370
rect 20778 24294 20886 24370
rect 0 24198 28 24246
rect 330 24040 438 24150
rect 810 24040 918 24150
rect 1578 24040 1686 24150
rect 2058 24040 2166 24150
rect 2826 24040 2934 24150
rect 3306 24040 3414 24150
rect 4074 24040 4182 24150
rect 4554 24040 4662 24150
rect 5322 24040 5430 24150
rect 5802 24040 5910 24150
rect 6570 24040 6678 24150
rect 7050 24040 7158 24150
rect 7818 24040 7926 24150
rect 8298 24040 8406 24150
rect 9066 24040 9174 24150
rect 9546 24040 9654 24150
rect 10314 24040 10422 24150
rect 10794 24040 10902 24150
rect 11562 24040 11670 24150
rect 12042 24040 12150 24150
rect 12810 24040 12918 24150
rect 13290 24040 13398 24150
rect 14058 24040 14166 24150
rect 14538 24040 14646 24150
rect 15306 24040 15414 24150
rect 15786 24040 15894 24150
rect 16554 24040 16662 24150
rect 17034 24040 17142 24150
rect 17802 24040 17910 24150
rect 18282 24040 18390 24150
rect 19050 24040 19158 24150
rect 19530 24040 19638 24150
rect 20298 24040 20406 24150
rect 20778 24040 20886 24150
rect 0 23944 28 23992
rect 330 23820 438 23896
rect 810 23820 918 23896
rect 1578 23820 1686 23896
rect 2058 23820 2166 23896
rect 2826 23820 2934 23896
rect 3306 23820 3414 23896
rect 4074 23820 4182 23896
rect 4554 23820 4662 23896
rect 5322 23820 5430 23896
rect 5802 23820 5910 23896
rect 6570 23820 6678 23896
rect 7050 23820 7158 23896
rect 7818 23820 7926 23896
rect 8298 23820 8406 23896
rect 9066 23820 9174 23896
rect 9546 23820 9654 23896
rect 10314 23820 10422 23896
rect 10794 23820 10902 23896
rect 11562 23820 11670 23896
rect 12042 23820 12150 23896
rect 12810 23820 12918 23896
rect 13290 23820 13398 23896
rect 14058 23820 14166 23896
rect 14538 23820 14646 23896
rect 15306 23820 15414 23896
rect 15786 23820 15894 23896
rect 16554 23820 16662 23896
rect 17034 23820 17142 23896
rect 17802 23820 17910 23896
rect 18282 23820 18390 23896
rect 19050 23820 19158 23896
rect 19530 23820 19638 23896
rect 20298 23820 20406 23896
rect 20778 23820 20886 23896
rect 0 23724 28 23772
rect 0 23628 28 23676
rect 330 23504 438 23580
rect 810 23504 918 23580
rect 1578 23504 1686 23580
rect 2058 23504 2166 23580
rect 2826 23504 2934 23580
rect 3306 23504 3414 23580
rect 4074 23504 4182 23580
rect 4554 23504 4662 23580
rect 5322 23504 5430 23580
rect 5802 23504 5910 23580
rect 6570 23504 6678 23580
rect 7050 23504 7158 23580
rect 7818 23504 7926 23580
rect 8298 23504 8406 23580
rect 9066 23504 9174 23580
rect 9546 23504 9654 23580
rect 10314 23504 10422 23580
rect 10794 23504 10902 23580
rect 11562 23504 11670 23580
rect 12042 23504 12150 23580
rect 12810 23504 12918 23580
rect 13290 23504 13398 23580
rect 14058 23504 14166 23580
rect 14538 23504 14646 23580
rect 15306 23504 15414 23580
rect 15786 23504 15894 23580
rect 16554 23504 16662 23580
rect 17034 23504 17142 23580
rect 17802 23504 17910 23580
rect 18282 23504 18390 23580
rect 19050 23504 19158 23580
rect 19530 23504 19638 23580
rect 20298 23504 20406 23580
rect 20778 23504 20886 23580
rect 0 23408 28 23456
rect 330 23250 438 23360
rect 810 23250 918 23360
rect 1578 23250 1686 23360
rect 2058 23250 2166 23360
rect 2826 23250 2934 23360
rect 3306 23250 3414 23360
rect 4074 23250 4182 23360
rect 4554 23250 4662 23360
rect 5322 23250 5430 23360
rect 5802 23250 5910 23360
rect 6570 23250 6678 23360
rect 7050 23250 7158 23360
rect 7818 23250 7926 23360
rect 8298 23250 8406 23360
rect 9066 23250 9174 23360
rect 9546 23250 9654 23360
rect 10314 23250 10422 23360
rect 10794 23250 10902 23360
rect 11562 23250 11670 23360
rect 12042 23250 12150 23360
rect 12810 23250 12918 23360
rect 13290 23250 13398 23360
rect 14058 23250 14166 23360
rect 14538 23250 14646 23360
rect 15306 23250 15414 23360
rect 15786 23250 15894 23360
rect 16554 23250 16662 23360
rect 17034 23250 17142 23360
rect 17802 23250 17910 23360
rect 18282 23250 18390 23360
rect 19050 23250 19158 23360
rect 19530 23250 19638 23360
rect 20298 23250 20406 23360
rect 20778 23250 20886 23360
rect 0 23154 28 23202
rect 330 23030 438 23106
rect 810 23030 918 23106
rect 1578 23030 1686 23106
rect 2058 23030 2166 23106
rect 2826 23030 2934 23106
rect 3306 23030 3414 23106
rect 4074 23030 4182 23106
rect 4554 23030 4662 23106
rect 5322 23030 5430 23106
rect 5802 23030 5910 23106
rect 6570 23030 6678 23106
rect 7050 23030 7158 23106
rect 7818 23030 7926 23106
rect 8298 23030 8406 23106
rect 9066 23030 9174 23106
rect 9546 23030 9654 23106
rect 10314 23030 10422 23106
rect 10794 23030 10902 23106
rect 11562 23030 11670 23106
rect 12042 23030 12150 23106
rect 12810 23030 12918 23106
rect 13290 23030 13398 23106
rect 14058 23030 14166 23106
rect 14538 23030 14646 23106
rect 15306 23030 15414 23106
rect 15786 23030 15894 23106
rect 16554 23030 16662 23106
rect 17034 23030 17142 23106
rect 17802 23030 17910 23106
rect 18282 23030 18390 23106
rect 19050 23030 19158 23106
rect 19530 23030 19638 23106
rect 20298 23030 20406 23106
rect 20778 23030 20886 23106
rect 0 22934 28 22982
rect 0 22838 28 22886
rect 330 22714 438 22790
rect 810 22714 918 22790
rect 1578 22714 1686 22790
rect 2058 22714 2166 22790
rect 2826 22714 2934 22790
rect 3306 22714 3414 22790
rect 4074 22714 4182 22790
rect 4554 22714 4662 22790
rect 5322 22714 5430 22790
rect 5802 22714 5910 22790
rect 6570 22714 6678 22790
rect 7050 22714 7158 22790
rect 7818 22714 7926 22790
rect 8298 22714 8406 22790
rect 9066 22714 9174 22790
rect 9546 22714 9654 22790
rect 10314 22714 10422 22790
rect 10794 22714 10902 22790
rect 11562 22714 11670 22790
rect 12042 22714 12150 22790
rect 12810 22714 12918 22790
rect 13290 22714 13398 22790
rect 14058 22714 14166 22790
rect 14538 22714 14646 22790
rect 15306 22714 15414 22790
rect 15786 22714 15894 22790
rect 16554 22714 16662 22790
rect 17034 22714 17142 22790
rect 17802 22714 17910 22790
rect 18282 22714 18390 22790
rect 19050 22714 19158 22790
rect 19530 22714 19638 22790
rect 20298 22714 20406 22790
rect 20778 22714 20886 22790
rect 0 22618 28 22666
rect 330 22460 438 22570
rect 810 22460 918 22570
rect 1578 22460 1686 22570
rect 2058 22460 2166 22570
rect 2826 22460 2934 22570
rect 3306 22460 3414 22570
rect 4074 22460 4182 22570
rect 4554 22460 4662 22570
rect 5322 22460 5430 22570
rect 5802 22460 5910 22570
rect 6570 22460 6678 22570
rect 7050 22460 7158 22570
rect 7818 22460 7926 22570
rect 8298 22460 8406 22570
rect 9066 22460 9174 22570
rect 9546 22460 9654 22570
rect 10314 22460 10422 22570
rect 10794 22460 10902 22570
rect 11562 22460 11670 22570
rect 12042 22460 12150 22570
rect 12810 22460 12918 22570
rect 13290 22460 13398 22570
rect 14058 22460 14166 22570
rect 14538 22460 14646 22570
rect 15306 22460 15414 22570
rect 15786 22460 15894 22570
rect 16554 22460 16662 22570
rect 17034 22460 17142 22570
rect 17802 22460 17910 22570
rect 18282 22460 18390 22570
rect 19050 22460 19158 22570
rect 19530 22460 19638 22570
rect 20298 22460 20406 22570
rect 20778 22460 20886 22570
rect 0 22364 28 22412
rect 330 22240 438 22316
rect 810 22240 918 22316
rect 1578 22240 1686 22316
rect 2058 22240 2166 22316
rect 2826 22240 2934 22316
rect 3306 22240 3414 22316
rect 4074 22240 4182 22316
rect 4554 22240 4662 22316
rect 5322 22240 5430 22316
rect 5802 22240 5910 22316
rect 6570 22240 6678 22316
rect 7050 22240 7158 22316
rect 7818 22240 7926 22316
rect 8298 22240 8406 22316
rect 9066 22240 9174 22316
rect 9546 22240 9654 22316
rect 10314 22240 10422 22316
rect 10794 22240 10902 22316
rect 11562 22240 11670 22316
rect 12042 22240 12150 22316
rect 12810 22240 12918 22316
rect 13290 22240 13398 22316
rect 14058 22240 14166 22316
rect 14538 22240 14646 22316
rect 15306 22240 15414 22316
rect 15786 22240 15894 22316
rect 16554 22240 16662 22316
rect 17034 22240 17142 22316
rect 17802 22240 17910 22316
rect 18282 22240 18390 22316
rect 19050 22240 19158 22316
rect 19530 22240 19638 22316
rect 20298 22240 20406 22316
rect 20778 22240 20886 22316
rect 0 22144 28 22192
rect 0 22048 28 22096
rect 330 21924 438 22000
rect 810 21924 918 22000
rect 1578 21924 1686 22000
rect 2058 21924 2166 22000
rect 2826 21924 2934 22000
rect 3306 21924 3414 22000
rect 4074 21924 4182 22000
rect 4554 21924 4662 22000
rect 5322 21924 5430 22000
rect 5802 21924 5910 22000
rect 6570 21924 6678 22000
rect 7050 21924 7158 22000
rect 7818 21924 7926 22000
rect 8298 21924 8406 22000
rect 9066 21924 9174 22000
rect 9546 21924 9654 22000
rect 10314 21924 10422 22000
rect 10794 21924 10902 22000
rect 11562 21924 11670 22000
rect 12042 21924 12150 22000
rect 12810 21924 12918 22000
rect 13290 21924 13398 22000
rect 14058 21924 14166 22000
rect 14538 21924 14646 22000
rect 15306 21924 15414 22000
rect 15786 21924 15894 22000
rect 16554 21924 16662 22000
rect 17034 21924 17142 22000
rect 17802 21924 17910 22000
rect 18282 21924 18390 22000
rect 19050 21924 19158 22000
rect 19530 21924 19638 22000
rect 20298 21924 20406 22000
rect 20778 21924 20886 22000
rect 0 21828 28 21876
rect 330 21670 438 21780
rect 810 21670 918 21780
rect 1578 21670 1686 21780
rect 2058 21670 2166 21780
rect 2826 21670 2934 21780
rect 3306 21670 3414 21780
rect 4074 21670 4182 21780
rect 4554 21670 4662 21780
rect 5322 21670 5430 21780
rect 5802 21670 5910 21780
rect 6570 21670 6678 21780
rect 7050 21670 7158 21780
rect 7818 21670 7926 21780
rect 8298 21670 8406 21780
rect 9066 21670 9174 21780
rect 9546 21670 9654 21780
rect 10314 21670 10422 21780
rect 10794 21670 10902 21780
rect 11562 21670 11670 21780
rect 12042 21670 12150 21780
rect 12810 21670 12918 21780
rect 13290 21670 13398 21780
rect 14058 21670 14166 21780
rect 14538 21670 14646 21780
rect 15306 21670 15414 21780
rect 15786 21670 15894 21780
rect 16554 21670 16662 21780
rect 17034 21670 17142 21780
rect 17802 21670 17910 21780
rect 18282 21670 18390 21780
rect 19050 21670 19158 21780
rect 19530 21670 19638 21780
rect 20298 21670 20406 21780
rect 20778 21670 20886 21780
rect 0 21574 28 21622
rect 330 21450 438 21526
rect 810 21450 918 21526
rect 1578 21450 1686 21526
rect 2058 21450 2166 21526
rect 2826 21450 2934 21526
rect 3306 21450 3414 21526
rect 4074 21450 4182 21526
rect 4554 21450 4662 21526
rect 5322 21450 5430 21526
rect 5802 21450 5910 21526
rect 6570 21450 6678 21526
rect 7050 21450 7158 21526
rect 7818 21450 7926 21526
rect 8298 21450 8406 21526
rect 9066 21450 9174 21526
rect 9546 21450 9654 21526
rect 10314 21450 10422 21526
rect 10794 21450 10902 21526
rect 11562 21450 11670 21526
rect 12042 21450 12150 21526
rect 12810 21450 12918 21526
rect 13290 21450 13398 21526
rect 14058 21450 14166 21526
rect 14538 21450 14646 21526
rect 15306 21450 15414 21526
rect 15786 21450 15894 21526
rect 16554 21450 16662 21526
rect 17034 21450 17142 21526
rect 17802 21450 17910 21526
rect 18282 21450 18390 21526
rect 19050 21450 19158 21526
rect 19530 21450 19638 21526
rect 20298 21450 20406 21526
rect 20778 21450 20886 21526
rect 0 21354 28 21402
rect 0 21258 28 21306
rect 330 21134 438 21210
rect 810 21134 918 21210
rect 1578 21134 1686 21210
rect 2058 21134 2166 21210
rect 2826 21134 2934 21210
rect 3306 21134 3414 21210
rect 4074 21134 4182 21210
rect 4554 21134 4662 21210
rect 5322 21134 5430 21210
rect 5802 21134 5910 21210
rect 6570 21134 6678 21210
rect 7050 21134 7158 21210
rect 7818 21134 7926 21210
rect 8298 21134 8406 21210
rect 9066 21134 9174 21210
rect 9546 21134 9654 21210
rect 10314 21134 10422 21210
rect 10794 21134 10902 21210
rect 11562 21134 11670 21210
rect 12042 21134 12150 21210
rect 12810 21134 12918 21210
rect 13290 21134 13398 21210
rect 14058 21134 14166 21210
rect 14538 21134 14646 21210
rect 15306 21134 15414 21210
rect 15786 21134 15894 21210
rect 16554 21134 16662 21210
rect 17034 21134 17142 21210
rect 17802 21134 17910 21210
rect 18282 21134 18390 21210
rect 19050 21134 19158 21210
rect 19530 21134 19638 21210
rect 20298 21134 20406 21210
rect 20778 21134 20886 21210
rect 0 21038 28 21086
rect 330 20880 438 20990
rect 810 20880 918 20990
rect 1578 20880 1686 20990
rect 2058 20880 2166 20990
rect 2826 20880 2934 20990
rect 3306 20880 3414 20990
rect 4074 20880 4182 20990
rect 4554 20880 4662 20990
rect 5322 20880 5430 20990
rect 5802 20880 5910 20990
rect 6570 20880 6678 20990
rect 7050 20880 7158 20990
rect 7818 20880 7926 20990
rect 8298 20880 8406 20990
rect 9066 20880 9174 20990
rect 9546 20880 9654 20990
rect 10314 20880 10422 20990
rect 10794 20880 10902 20990
rect 11562 20880 11670 20990
rect 12042 20880 12150 20990
rect 12810 20880 12918 20990
rect 13290 20880 13398 20990
rect 14058 20880 14166 20990
rect 14538 20880 14646 20990
rect 15306 20880 15414 20990
rect 15786 20880 15894 20990
rect 16554 20880 16662 20990
rect 17034 20880 17142 20990
rect 17802 20880 17910 20990
rect 18282 20880 18390 20990
rect 19050 20880 19158 20990
rect 19530 20880 19638 20990
rect 20298 20880 20406 20990
rect 20778 20880 20886 20990
rect 0 20784 28 20832
rect 330 20660 438 20736
rect 810 20660 918 20736
rect 1578 20660 1686 20736
rect 2058 20660 2166 20736
rect 2826 20660 2934 20736
rect 3306 20660 3414 20736
rect 4074 20660 4182 20736
rect 4554 20660 4662 20736
rect 5322 20660 5430 20736
rect 5802 20660 5910 20736
rect 6570 20660 6678 20736
rect 7050 20660 7158 20736
rect 7818 20660 7926 20736
rect 8298 20660 8406 20736
rect 9066 20660 9174 20736
rect 9546 20660 9654 20736
rect 10314 20660 10422 20736
rect 10794 20660 10902 20736
rect 11562 20660 11670 20736
rect 12042 20660 12150 20736
rect 12810 20660 12918 20736
rect 13290 20660 13398 20736
rect 14058 20660 14166 20736
rect 14538 20660 14646 20736
rect 15306 20660 15414 20736
rect 15786 20660 15894 20736
rect 16554 20660 16662 20736
rect 17034 20660 17142 20736
rect 17802 20660 17910 20736
rect 18282 20660 18390 20736
rect 19050 20660 19158 20736
rect 19530 20660 19638 20736
rect 20298 20660 20406 20736
rect 20778 20660 20886 20736
rect 0 20564 28 20612
rect 0 20468 28 20516
rect 330 20344 438 20420
rect 810 20344 918 20420
rect 1578 20344 1686 20420
rect 2058 20344 2166 20420
rect 2826 20344 2934 20420
rect 3306 20344 3414 20420
rect 4074 20344 4182 20420
rect 4554 20344 4662 20420
rect 5322 20344 5430 20420
rect 5802 20344 5910 20420
rect 6570 20344 6678 20420
rect 7050 20344 7158 20420
rect 7818 20344 7926 20420
rect 8298 20344 8406 20420
rect 9066 20344 9174 20420
rect 9546 20344 9654 20420
rect 10314 20344 10422 20420
rect 10794 20344 10902 20420
rect 11562 20344 11670 20420
rect 12042 20344 12150 20420
rect 12810 20344 12918 20420
rect 13290 20344 13398 20420
rect 14058 20344 14166 20420
rect 14538 20344 14646 20420
rect 15306 20344 15414 20420
rect 15786 20344 15894 20420
rect 16554 20344 16662 20420
rect 17034 20344 17142 20420
rect 17802 20344 17910 20420
rect 18282 20344 18390 20420
rect 19050 20344 19158 20420
rect 19530 20344 19638 20420
rect 20298 20344 20406 20420
rect 20778 20344 20886 20420
rect 0 20248 28 20296
rect 330 20090 438 20200
rect 810 20090 918 20200
rect 1578 20090 1686 20200
rect 2058 20090 2166 20200
rect 2826 20090 2934 20200
rect 3306 20090 3414 20200
rect 4074 20090 4182 20200
rect 4554 20090 4662 20200
rect 5322 20090 5430 20200
rect 5802 20090 5910 20200
rect 6570 20090 6678 20200
rect 7050 20090 7158 20200
rect 7818 20090 7926 20200
rect 8298 20090 8406 20200
rect 9066 20090 9174 20200
rect 9546 20090 9654 20200
rect 10314 20090 10422 20200
rect 10794 20090 10902 20200
rect 11562 20090 11670 20200
rect 12042 20090 12150 20200
rect 12810 20090 12918 20200
rect 13290 20090 13398 20200
rect 14058 20090 14166 20200
rect 14538 20090 14646 20200
rect 15306 20090 15414 20200
rect 15786 20090 15894 20200
rect 16554 20090 16662 20200
rect 17034 20090 17142 20200
rect 17802 20090 17910 20200
rect 18282 20090 18390 20200
rect 19050 20090 19158 20200
rect 19530 20090 19638 20200
rect 20298 20090 20406 20200
rect 20778 20090 20886 20200
rect 0 19994 28 20042
rect 330 19870 438 19946
rect 810 19870 918 19946
rect 1578 19870 1686 19946
rect 2058 19870 2166 19946
rect 2826 19870 2934 19946
rect 3306 19870 3414 19946
rect 4074 19870 4182 19946
rect 4554 19870 4662 19946
rect 5322 19870 5430 19946
rect 5802 19870 5910 19946
rect 6570 19870 6678 19946
rect 7050 19870 7158 19946
rect 7818 19870 7926 19946
rect 8298 19870 8406 19946
rect 9066 19870 9174 19946
rect 9546 19870 9654 19946
rect 10314 19870 10422 19946
rect 10794 19870 10902 19946
rect 11562 19870 11670 19946
rect 12042 19870 12150 19946
rect 12810 19870 12918 19946
rect 13290 19870 13398 19946
rect 14058 19870 14166 19946
rect 14538 19870 14646 19946
rect 15306 19870 15414 19946
rect 15786 19870 15894 19946
rect 16554 19870 16662 19946
rect 17034 19870 17142 19946
rect 17802 19870 17910 19946
rect 18282 19870 18390 19946
rect 19050 19870 19158 19946
rect 19530 19870 19638 19946
rect 20298 19870 20406 19946
rect 20778 19870 20886 19946
rect 0 19774 28 19822
rect 0 19678 28 19726
rect 330 19554 438 19630
rect 810 19554 918 19630
rect 1578 19554 1686 19630
rect 2058 19554 2166 19630
rect 2826 19554 2934 19630
rect 3306 19554 3414 19630
rect 4074 19554 4182 19630
rect 4554 19554 4662 19630
rect 5322 19554 5430 19630
rect 5802 19554 5910 19630
rect 6570 19554 6678 19630
rect 7050 19554 7158 19630
rect 7818 19554 7926 19630
rect 8298 19554 8406 19630
rect 9066 19554 9174 19630
rect 9546 19554 9654 19630
rect 10314 19554 10422 19630
rect 10794 19554 10902 19630
rect 11562 19554 11670 19630
rect 12042 19554 12150 19630
rect 12810 19554 12918 19630
rect 13290 19554 13398 19630
rect 14058 19554 14166 19630
rect 14538 19554 14646 19630
rect 15306 19554 15414 19630
rect 15786 19554 15894 19630
rect 16554 19554 16662 19630
rect 17034 19554 17142 19630
rect 17802 19554 17910 19630
rect 18282 19554 18390 19630
rect 19050 19554 19158 19630
rect 19530 19554 19638 19630
rect 20298 19554 20406 19630
rect 20778 19554 20886 19630
rect 0 19458 28 19506
rect 330 19300 438 19410
rect 810 19300 918 19410
rect 1578 19300 1686 19410
rect 2058 19300 2166 19410
rect 2826 19300 2934 19410
rect 3306 19300 3414 19410
rect 4074 19300 4182 19410
rect 4554 19300 4662 19410
rect 5322 19300 5430 19410
rect 5802 19300 5910 19410
rect 6570 19300 6678 19410
rect 7050 19300 7158 19410
rect 7818 19300 7926 19410
rect 8298 19300 8406 19410
rect 9066 19300 9174 19410
rect 9546 19300 9654 19410
rect 10314 19300 10422 19410
rect 10794 19300 10902 19410
rect 11562 19300 11670 19410
rect 12042 19300 12150 19410
rect 12810 19300 12918 19410
rect 13290 19300 13398 19410
rect 14058 19300 14166 19410
rect 14538 19300 14646 19410
rect 15306 19300 15414 19410
rect 15786 19300 15894 19410
rect 16554 19300 16662 19410
rect 17034 19300 17142 19410
rect 17802 19300 17910 19410
rect 18282 19300 18390 19410
rect 19050 19300 19158 19410
rect 19530 19300 19638 19410
rect 20298 19300 20406 19410
rect 20778 19300 20886 19410
rect 0 19204 28 19252
rect 330 19080 438 19156
rect 810 19080 918 19156
rect 1578 19080 1686 19156
rect 2058 19080 2166 19156
rect 2826 19080 2934 19156
rect 3306 19080 3414 19156
rect 4074 19080 4182 19156
rect 4554 19080 4662 19156
rect 5322 19080 5430 19156
rect 5802 19080 5910 19156
rect 6570 19080 6678 19156
rect 7050 19080 7158 19156
rect 7818 19080 7926 19156
rect 8298 19080 8406 19156
rect 9066 19080 9174 19156
rect 9546 19080 9654 19156
rect 10314 19080 10422 19156
rect 10794 19080 10902 19156
rect 11562 19080 11670 19156
rect 12042 19080 12150 19156
rect 12810 19080 12918 19156
rect 13290 19080 13398 19156
rect 14058 19080 14166 19156
rect 14538 19080 14646 19156
rect 15306 19080 15414 19156
rect 15786 19080 15894 19156
rect 16554 19080 16662 19156
rect 17034 19080 17142 19156
rect 17802 19080 17910 19156
rect 18282 19080 18390 19156
rect 19050 19080 19158 19156
rect 19530 19080 19638 19156
rect 20298 19080 20406 19156
rect 20778 19080 20886 19156
rect 0 18984 28 19032
rect 0 18888 28 18936
rect 330 18764 438 18840
rect 810 18764 918 18840
rect 1578 18764 1686 18840
rect 2058 18764 2166 18840
rect 2826 18764 2934 18840
rect 3306 18764 3414 18840
rect 4074 18764 4182 18840
rect 4554 18764 4662 18840
rect 5322 18764 5430 18840
rect 5802 18764 5910 18840
rect 6570 18764 6678 18840
rect 7050 18764 7158 18840
rect 7818 18764 7926 18840
rect 8298 18764 8406 18840
rect 9066 18764 9174 18840
rect 9546 18764 9654 18840
rect 10314 18764 10422 18840
rect 10794 18764 10902 18840
rect 11562 18764 11670 18840
rect 12042 18764 12150 18840
rect 12810 18764 12918 18840
rect 13290 18764 13398 18840
rect 14058 18764 14166 18840
rect 14538 18764 14646 18840
rect 15306 18764 15414 18840
rect 15786 18764 15894 18840
rect 16554 18764 16662 18840
rect 17034 18764 17142 18840
rect 17802 18764 17910 18840
rect 18282 18764 18390 18840
rect 19050 18764 19158 18840
rect 19530 18764 19638 18840
rect 20298 18764 20406 18840
rect 20778 18764 20886 18840
rect 0 18668 28 18716
rect 330 18510 438 18620
rect 810 18510 918 18620
rect 1578 18510 1686 18620
rect 2058 18510 2166 18620
rect 2826 18510 2934 18620
rect 3306 18510 3414 18620
rect 4074 18510 4182 18620
rect 4554 18510 4662 18620
rect 5322 18510 5430 18620
rect 5802 18510 5910 18620
rect 6570 18510 6678 18620
rect 7050 18510 7158 18620
rect 7818 18510 7926 18620
rect 8298 18510 8406 18620
rect 9066 18510 9174 18620
rect 9546 18510 9654 18620
rect 10314 18510 10422 18620
rect 10794 18510 10902 18620
rect 11562 18510 11670 18620
rect 12042 18510 12150 18620
rect 12810 18510 12918 18620
rect 13290 18510 13398 18620
rect 14058 18510 14166 18620
rect 14538 18510 14646 18620
rect 15306 18510 15414 18620
rect 15786 18510 15894 18620
rect 16554 18510 16662 18620
rect 17034 18510 17142 18620
rect 17802 18510 17910 18620
rect 18282 18510 18390 18620
rect 19050 18510 19158 18620
rect 19530 18510 19638 18620
rect 20298 18510 20406 18620
rect 20778 18510 20886 18620
rect 0 18414 28 18462
rect 330 18290 438 18366
rect 810 18290 918 18366
rect 1578 18290 1686 18366
rect 2058 18290 2166 18366
rect 2826 18290 2934 18366
rect 3306 18290 3414 18366
rect 4074 18290 4182 18366
rect 4554 18290 4662 18366
rect 5322 18290 5430 18366
rect 5802 18290 5910 18366
rect 6570 18290 6678 18366
rect 7050 18290 7158 18366
rect 7818 18290 7926 18366
rect 8298 18290 8406 18366
rect 9066 18290 9174 18366
rect 9546 18290 9654 18366
rect 10314 18290 10422 18366
rect 10794 18290 10902 18366
rect 11562 18290 11670 18366
rect 12042 18290 12150 18366
rect 12810 18290 12918 18366
rect 13290 18290 13398 18366
rect 14058 18290 14166 18366
rect 14538 18290 14646 18366
rect 15306 18290 15414 18366
rect 15786 18290 15894 18366
rect 16554 18290 16662 18366
rect 17034 18290 17142 18366
rect 17802 18290 17910 18366
rect 18282 18290 18390 18366
rect 19050 18290 19158 18366
rect 19530 18290 19638 18366
rect 20298 18290 20406 18366
rect 20778 18290 20886 18366
rect 0 18194 28 18242
rect 0 18098 28 18146
rect 330 17974 438 18050
rect 810 17974 918 18050
rect 1578 17974 1686 18050
rect 2058 17974 2166 18050
rect 2826 17974 2934 18050
rect 3306 17974 3414 18050
rect 4074 17974 4182 18050
rect 4554 17974 4662 18050
rect 5322 17974 5430 18050
rect 5802 17974 5910 18050
rect 6570 17974 6678 18050
rect 7050 17974 7158 18050
rect 7818 17974 7926 18050
rect 8298 17974 8406 18050
rect 9066 17974 9174 18050
rect 9546 17974 9654 18050
rect 10314 17974 10422 18050
rect 10794 17974 10902 18050
rect 11562 17974 11670 18050
rect 12042 17974 12150 18050
rect 12810 17974 12918 18050
rect 13290 17974 13398 18050
rect 14058 17974 14166 18050
rect 14538 17974 14646 18050
rect 15306 17974 15414 18050
rect 15786 17974 15894 18050
rect 16554 17974 16662 18050
rect 17034 17974 17142 18050
rect 17802 17974 17910 18050
rect 18282 17974 18390 18050
rect 19050 17974 19158 18050
rect 19530 17974 19638 18050
rect 20298 17974 20406 18050
rect 20778 17974 20886 18050
rect 0 17878 28 17926
rect 330 17720 438 17830
rect 810 17720 918 17830
rect 1578 17720 1686 17830
rect 2058 17720 2166 17830
rect 2826 17720 2934 17830
rect 3306 17720 3414 17830
rect 4074 17720 4182 17830
rect 4554 17720 4662 17830
rect 5322 17720 5430 17830
rect 5802 17720 5910 17830
rect 6570 17720 6678 17830
rect 7050 17720 7158 17830
rect 7818 17720 7926 17830
rect 8298 17720 8406 17830
rect 9066 17720 9174 17830
rect 9546 17720 9654 17830
rect 10314 17720 10422 17830
rect 10794 17720 10902 17830
rect 11562 17720 11670 17830
rect 12042 17720 12150 17830
rect 12810 17720 12918 17830
rect 13290 17720 13398 17830
rect 14058 17720 14166 17830
rect 14538 17720 14646 17830
rect 15306 17720 15414 17830
rect 15786 17720 15894 17830
rect 16554 17720 16662 17830
rect 17034 17720 17142 17830
rect 17802 17720 17910 17830
rect 18282 17720 18390 17830
rect 19050 17720 19158 17830
rect 19530 17720 19638 17830
rect 20298 17720 20406 17830
rect 20778 17720 20886 17830
rect 0 17624 28 17672
rect 330 17500 438 17576
rect 810 17500 918 17576
rect 1578 17500 1686 17576
rect 2058 17500 2166 17576
rect 2826 17500 2934 17576
rect 3306 17500 3414 17576
rect 4074 17500 4182 17576
rect 4554 17500 4662 17576
rect 5322 17500 5430 17576
rect 5802 17500 5910 17576
rect 6570 17500 6678 17576
rect 7050 17500 7158 17576
rect 7818 17500 7926 17576
rect 8298 17500 8406 17576
rect 9066 17500 9174 17576
rect 9546 17500 9654 17576
rect 10314 17500 10422 17576
rect 10794 17500 10902 17576
rect 11562 17500 11670 17576
rect 12042 17500 12150 17576
rect 12810 17500 12918 17576
rect 13290 17500 13398 17576
rect 14058 17500 14166 17576
rect 14538 17500 14646 17576
rect 15306 17500 15414 17576
rect 15786 17500 15894 17576
rect 16554 17500 16662 17576
rect 17034 17500 17142 17576
rect 17802 17500 17910 17576
rect 18282 17500 18390 17576
rect 19050 17500 19158 17576
rect 19530 17500 19638 17576
rect 20298 17500 20406 17576
rect 20778 17500 20886 17576
rect 0 17404 28 17452
rect 0 17308 28 17356
rect 330 17184 438 17260
rect 810 17184 918 17260
rect 1578 17184 1686 17260
rect 2058 17184 2166 17260
rect 2826 17184 2934 17260
rect 3306 17184 3414 17260
rect 4074 17184 4182 17260
rect 4554 17184 4662 17260
rect 5322 17184 5430 17260
rect 5802 17184 5910 17260
rect 6570 17184 6678 17260
rect 7050 17184 7158 17260
rect 7818 17184 7926 17260
rect 8298 17184 8406 17260
rect 9066 17184 9174 17260
rect 9546 17184 9654 17260
rect 10314 17184 10422 17260
rect 10794 17184 10902 17260
rect 11562 17184 11670 17260
rect 12042 17184 12150 17260
rect 12810 17184 12918 17260
rect 13290 17184 13398 17260
rect 14058 17184 14166 17260
rect 14538 17184 14646 17260
rect 15306 17184 15414 17260
rect 15786 17184 15894 17260
rect 16554 17184 16662 17260
rect 17034 17184 17142 17260
rect 17802 17184 17910 17260
rect 18282 17184 18390 17260
rect 19050 17184 19158 17260
rect 19530 17184 19638 17260
rect 20298 17184 20406 17260
rect 20778 17184 20886 17260
rect 0 17088 28 17136
rect 330 16930 438 17040
rect 810 16930 918 17040
rect 1578 16930 1686 17040
rect 2058 16930 2166 17040
rect 2826 16930 2934 17040
rect 3306 16930 3414 17040
rect 4074 16930 4182 17040
rect 4554 16930 4662 17040
rect 5322 16930 5430 17040
rect 5802 16930 5910 17040
rect 6570 16930 6678 17040
rect 7050 16930 7158 17040
rect 7818 16930 7926 17040
rect 8298 16930 8406 17040
rect 9066 16930 9174 17040
rect 9546 16930 9654 17040
rect 10314 16930 10422 17040
rect 10794 16930 10902 17040
rect 11562 16930 11670 17040
rect 12042 16930 12150 17040
rect 12810 16930 12918 17040
rect 13290 16930 13398 17040
rect 14058 16930 14166 17040
rect 14538 16930 14646 17040
rect 15306 16930 15414 17040
rect 15786 16930 15894 17040
rect 16554 16930 16662 17040
rect 17034 16930 17142 17040
rect 17802 16930 17910 17040
rect 18282 16930 18390 17040
rect 19050 16930 19158 17040
rect 19530 16930 19638 17040
rect 20298 16930 20406 17040
rect 20778 16930 20886 17040
rect 0 16834 28 16882
rect 330 16710 438 16786
rect 810 16710 918 16786
rect 1578 16710 1686 16786
rect 2058 16710 2166 16786
rect 2826 16710 2934 16786
rect 3306 16710 3414 16786
rect 4074 16710 4182 16786
rect 4554 16710 4662 16786
rect 5322 16710 5430 16786
rect 5802 16710 5910 16786
rect 6570 16710 6678 16786
rect 7050 16710 7158 16786
rect 7818 16710 7926 16786
rect 8298 16710 8406 16786
rect 9066 16710 9174 16786
rect 9546 16710 9654 16786
rect 10314 16710 10422 16786
rect 10794 16710 10902 16786
rect 11562 16710 11670 16786
rect 12042 16710 12150 16786
rect 12810 16710 12918 16786
rect 13290 16710 13398 16786
rect 14058 16710 14166 16786
rect 14538 16710 14646 16786
rect 15306 16710 15414 16786
rect 15786 16710 15894 16786
rect 16554 16710 16662 16786
rect 17034 16710 17142 16786
rect 17802 16710 17910 16786
rect 18282 16710 18390 16786
rect 19050 16710 19158 16786
rect 19530 16710 19638 16786
rect 20298 16710 20406 16786
rect 20778 16710 20886 16786
rect 0 16614 28 16662
rect 0 16518 28 16566
rect 330 16394 438 16470
rect 810 16394 918 16470
rect 1578 16394 1686 16470
rect 2058 16394 2166 16470
rect 2826 16394 2934 16470
rect 3306 16394 3414 16470
rect 4074 16394 4182 16470
rect 4554 16394 4662 16470
rect 5322 16394 5430 16470
rect 5802 16394 5910 16470
rect 6570 16394 6678 16470
rect 7050 16394 7158 16470
rect 7818 16394 7926 16470
rect 8298 16394 8406 16470
rect 9066 16394 9174 16470
rect 9546 16394 9654 16470
rect 10314 16394 10422 16470
rect 10794 16394 10902 16470
rect 11562 16394 11670 16470
rect 12042 16394 12150 16470
rect 12810 16394 12918 16470
rect 13290 16394 13398 16470
rect 14058 16394 14166 16470
rect 14538 16394 14646 16470
rect 15306 16394 15414 16470
rect 15786 16394 15894 16470
rect 16554 16394 16662 16470
rect 17034 16394 17142 16470
rect 17802 16394 17910 16470
rect 18282 16394 18390 16470
rect 19050 16394 19158 16470
rect 19530 16394 19638 16470
rect 20298 16394 20406 16470
rect 20778 16394 20886 16470
rect 0 16298 28 16346
rect 330 16140 438 16250
rect 810 16140 918 16250
rect 1578 16140 1686 16250
rect 2058 16140 2166 16250
rect 2826 16140 2934 16250
rect 3306 16140 3414 16250
rect 4074 16140 4182 16250
rect 4554 16140 4662 16250
rect 5322 16140 5430 16250
rect 5802 16140 5910 16250
rect 6570 16140 6678 16250
rect 7050 16140 7158 16250
rect 7818 16140 7926 16250
rect 8298 16140 8406 16250
rect 9066 16140 9174 16250
rect 9546 16140 9654 16250
rect 10314 16140 10422 16250
rect 10794 16140 10902 16250
rect 11562 16140 11670 16250
rect 12042 16140 12150 16250
rect 12810 16140 12918 16250
rect 13290 16140 13398 16250
rect 14058 16140 14166 16250
rect 14538 16140 14646 16250
rect 15306 16140 15414 16250
rect 15786 16140 15894 16250
rect 16554 16140 16662 16250
rect 17034 16140 17142 16250
rect 17802 16140 17910 16250
rect 18282 16140 18390 16250
rect 19050 16140 19158 16250
rect 19530 16140 19638 16250
rect 20298 16140 20406 16250
rect 20778 16140 20886 16250
rect 0 16044 28 16092
rect 330 15920 438 15996
rect 810 15920 918 15996
rect 1578 15920 1686 15996
rect 2058 15920 2166 15996
rect 2826 15920 2934 15996
rect 3306 15920 3414 15996
rect 4074 15920 4182 15996
rect 4554 15920 4662 15996
rect 5322 15920 5430 15996
rect 5802 15920 5910 15996
rect 6570 15920 6678 15996
rect 7050 15920 7158 15996
rect 7818 15920 7926 15996
rect 8298 15920 8406 15996
rect 9066 15920 9174 15996
rect 9546 15920 9654 15996
rect 10314 15920 10422 15996
rect 10794 15920 10902 15996
rect 11562 15920 11670 15996
rect 12042 15920 12150 15996
rect 12810 15920 12918 15996
rect 13290 15920 13398 15996
rect 14058 15920 14166 15996
rect 14538 15920 14646 15996
rect 15306 15920 15414 15996
rect 15786 15920 15894 15996
rect 16554 15920 16662 15996
rect 17034 15920 17142 15996
rect 17802 15920 17910 15996
rect 18282 15920 18390 15996
rect 19050 15920 19158 15996
rect 19530 15920 19638 15996
rect 20298 15920 20406 15996
rect 20778 15920 20886 15996
rect 0 15824 28 15872
rect 0 15728 28 15776
rect 330 15604 438 15680
rect 810 15604 918 15680
rect 1578 15604 1686 15680
rect 2058 15604 2166 15680
rect 2826 15604 2934 15680
rect 3306 15604 3414 15680
rect 4074 15604 4182 15680
rect 4554 15604 4662 15680
rect 5322 15604 5430 15680
rect 5802 15604 5910 15680
rect 6570 15604 6678 15680
rect 7050 15604 7158 15680
rect 7818 15604 7926 15680
rect 8298 15604 8406 15680
rect 9066 15604 9174 15680
rect 9546 15604 9654 15680
rect 10314 15604 10422 15680
rect 10794 15604 10902 15680
rect 11562 15604 11670 15680
rect 12042 15604 12150 15680
rect 12810 15604 12918 15680
rect 13290 15604 13398 15680
rect 14058 15604 14166 15680
rect 14538 15604 14646 15680
rect 15306 15604 15414 15680
rect 15786 15604 15894 15680
rect 16554 15604 16662 15680
rect 17034 15604 17142 15680
rect 17802 15604 17910 15680
rect 18282 15604 18390 15680
rect 19050 15604 19158 15680
rect 19530 15604 19638 15680
rect 20298 15604 20406 15680
rect 20778 15604 20886 15680
rect 0 15508 28 15556
rect 330 15350 438 15460
rect 810 15350 918 15460
rect 1578 15350 1686 15460
rect 2058 15350 2166 15460
rect 2826 15350 2934 15460
rect 3306 15350 3414 15460
rect 4074 15350 4182 15460
rect 4554 15350 4662 15460
rect 5322 15350 5430 15460
rect 5802 15350 5910 15460
rect 6570 15350 6678 15460
rect 7050 15350 7158 15460
rect 7818 15350 7926 15460
rect 8298 15350 8406 15460
rect 9066 15350 9174 15460
rect 9546 15350 9654 15460
rect 10314 15350 10422 15460
rect 10794 15350 10902 15460
rect 11562 15350 11670 15460
rect 12042 15350 12150 15460
rect 12810 15350 12918 15460
rect 13290 15350 13398 15460
rect 14058 15350 14166 15460
rect 14538 15350 14646 15460
rect 15306 15350 15414 15460
rect 15786 15350 15894 15460
rect 16554 15350 16662 15460
rect 17034 15350 17142 15460
rect 17802 15350 17910 15460
rect 18282 15350 18390 15460
rect 19050 15350 19158 15460
rect 19530 15350 19638 15460
rect 20298 15350 20406 15460
rect 20778 15350 20886 15460
rect 0 15254 28 15302
rect 330 15130 438 15206
rect 810 15130 918 15206
rect 1578 15130 1686 15206
rect 2058 15130 2166 15206
rect 2826 15130 2934 15206
rect 3306 15130 3414 15206
rect 4074 15130 4182 15206
rect 4554 15130 4662 15206
rect 5322 15130 5430 15206
rect 5802 15130 5910 15206
rect 6570 15130 6678 15206
rect 7050 15130 7158 15206
rect 7818 15130 7926 15206
rect 8298 15130 8406 15206
rect 9066 15130 9174 15206
rect 9546 15130 9654 15206
rect 10314 15130 10422 15206
rect 10794 15130 10902 15206
rect 11562 15130 11670 15206
rect 12042 15130 12150 15206
rect 12810 15130 12918 15206
rect 13290 15130 13398 15206
rect 14058 15130 14166 15206
rect 14538 15130 14646 15206
rect 15306 15130 15414 15206
rect 15786 15130 15894 15206
rect 16554 15130 16662 15206
rect 17034 15130 17142 15206
rect 17802 15130 17910 15206
rect 18282 15130 18390 15206
rect 19050 15130 19158 15206
rect 19530 15130 19638 15206
rect 20298 15130 20406 15206
rect 20778 15130 20886 15206
rect 0 15034 28 15082
rect 0 14938 28 14986
rect 330 14814 438 14890
rect 810 14814 918 14890
rect 1578 14814 1686 14890
rect 2058 14814 2166 14890
rect 2826 14814 2934 14890
rect 3306 14814 3414 14890
rect 4074 14814 4182 14890
rect 4554 14814 4662 14890
rect 5322 14814 5430 14890
rect 5802 14814 5910 14890
rect 6570 14814 6678 14890
rect 7050 14814 7158 14890
rect 7818 14814 7926 14890
rect 8298 14814 8406 14890
rect 9066 14814 9174 14890
rect 9546 14814 9654 14890
rect 10314 14814 10422 14890
rect 10794 14814 10902 14890
rect 11562 14814 11670 14890
rect 12042 14814 12150 14890
rect 12810 14814 12918 14890
rect 13290 14814 13398 14890
rect 14058 14814 14166 14890
rect 14538 14814 14646 14890
rect 15306 14814 15414 14890
rect 15786 14814 15894 14890
rect 16554 14814 16662 14890
rect 17034 14814 17142 14890
rect 17802 14814 17910 14890
rect 18282 14814 18390 14890
rect 19050 14814 19158 14890
rect 19530 14814 19638 14890
rect 20298 14814 20406 14890
rect 20778 14814 20886 14890
rect 0 14718 28 14766
rect 330 14560 438 14670
rect 810 14560 918 14670
rect 1578 14560 1686 14670
rect 2058 14560 2166 14670
rect 2826 14560 2934 14670
rect 3306 14560 3414 14670
rect 4074 14560 4182 14670
rect 4554 14560 4662 14670
rect 5322 14560 5430 14670
rect 5802 14560 5910 14670
rect 6570 14560 6678 14670
rect 7050 14560 7158 14670
rect 7818 14560 7926 14670
rect 8298 14560 8406 14670
rect 9066 14560 9174 14670
rect 9546 14560 9654 14670
rect 10314 14560 10422 14670
rect 10794 14560 10902 14670
rect 11562 14560 11670 14670
rect 12042 14560 12150 14670
rect 12810 14560 12918 14670
rect 13290 14560 13398 14670
rect 14058 14560 14166 14670
rect 14538 14560 14646 14670
rect 15306 14560 15414 14670
rect 15786 14560 15894 14670
rect 16554 14560 16662 14670
rect 17034 14560 17142 14670
rect 17802 14560 17910 14670
rect 18282 14560 18390 14670
rect 19050 14560 19158 14670
rect 19530 14560 19638 14670
rect 20298 14560 20406 14670
rect 20778 14560 20886 14670
rect 0 14464 28 14512
rect 330 14340 438 14416
rect 810 14340 918 14416
rect 1578 14340 1686 14416
rect 2058 14340 2166 14416
rect 2826 14340 2934 14416
rect 3306 14340 3414 14416
rect 4074 14340 4182 14416
rect 4554 14340 4662 14416
rect 5322 14340 5430 14416
rect 5802 14340 5910 14416
rect 6570 14340 6678 14416
rect 7050 14340 7158 14416
rect 7818 14340 7926 14416
rect 8298 14340 8406 14416
rect 9066 14340 9174 14416
rect 9546 14340 9654 14416
rect 10314 14340 10422 14416
rect 10794 14340 10902 14416
rect 11562 14340 11670 14416
rect 12042 14340 12150 14416
rect 12810 14340 12918 14416
rect 13290 14340 13398 14416
rect 14058 14340 14166 14416
rect 14538 14340 14646 14416
rect 15306 14340 15414 14416
rect 15786 14340 15894 14416
rect 16554 14340 16662 14416
rect 17034 14340 17142 14416
rect 17802 14340 17910 14416
rect 18282 14340 18390 14416
rect 19050 14340 19158 14416
rect 19530 14340 19638 14416
rect 20298 14340 20406 14416
rect 20778 14340 20886 14416
rect 0 14244 28 14292
rect 0 14148 28 14196
rect 330 14024 438 14100
rect 810 14024 918 14100
rect 1578 14024 1686 14100
rect 2058 14024 2166 14100
rect 2826 14024 2934 14100
rect 3306 14024 3414 14100
rect 4074 14024 4182 14100
rect 4554 14024 4662 14100
rect 5322 14024 5430 14100
rect 5802 14024 5910 14100
rect 6570 14024 6678 14100
rect 7050 14024 7158 14100
rect 7818 14024 7926 14100
rect 8298 14024 8406 14100
rect 9066 14024 9174 14100
rect 9546 14024 9654 14100
rect 10314 14024 10422 14100
rect 10794 14024 10902 14100
rect 11562 14024 11670 14100
rect 12042 14024 12150 14100
rect 12810 14024 12918 14100
rect 13290 14024 13398 14100
rect 14058 14024 14166 14100
rect 14538 14024 14646 14100
rect 15306 14024 15414 14100
rect 15786 14024 15894 14100
rect 16554 14024 16662 14100
rect 17034 14024 17142 14100
rect 17802 14024 17910 14100
rect 18282 14024 18390 14100
rect 19050 14024 19158 14100
rect 19530 14024 19638 14100
rect 20298 14024 20406 14100
rect 20778 14024 20886 14100
rect 0 13928 28 13976
rect 330 13770 438 13880
rect 810 13770 918 13880
rect 1578 13770 1686 13880
rect 2058 13770 2166 13880
rect 2826 13770 2934 13880
rect 3306 13770 3414 13880
rect 4074 13770 4182 13880
rect 4554 13770 4662 13880
rect 5322 13770 5430 13880
rect 5802 13770 5910 13880
rect 6570 13770 6678 13880
rect 7050 13770 7158 13880
rect 7818 13770 7926 13880
rect 8298 13770 8406 13880
rect 9066 13770 9174 13880
rect 9546 13770 9654 13880
rect 10314 13770 10422 13880
rect 10794 13770 10902 13880
rect 11562 13770 11670 13880
rect 12042 13770 12150 13880
rect 12810 13770 12918 13880
rect 13290 13770 13398 13880
rect 14058 13770 14166 13880
rect 14538 13770 14646 13880
rect 15306 13770 15414 13880
rect 15786 13770 15894 13880
rect 16554 13770 16662 13880
rect 17034 13770 17142 13880
rect 17802 13770 17910 13880
rect 18282 13770 18390 13880
rect 19050 13770 19158 13880
rect 19530 13770 19638 13880
rect 20298 13770 20406 13880
rect 20778 13770 20886 13880
rect 0 13674 28 13722
rect 330 13550 438 13626
rect 810 13550 918 13626
rect 1578 13550 1686 13626
rect 2058 13550 2166 13626
rect 2826 13550 2934 13626
rect 3306 13550 3414 13626
rect 4074 13550 4182 13626
rect 4554 13550 4662 13626
rect 5322 13550 5430 13626
rect 5802 13550 5910 13626
rect 6570 13550 6678 13626
rect 7050 13550 7158 13626
rect 7818 13550 7926 13626
rect 8298 13550 8406 13626
rect 9066 13550 9174 13626
rect 9546 13550 9654 13626
rect 10314 13550 10422 13626
rect 10794 13550 10902 13626
rect 11562 13550 11670 13626
rect 12042 13550 12150 13626
rect 12810 13550 12918 13626
rect 13290 13550 13398 13626
rect 14058 13550 14166 13626
rect 14538 13550 14646 13626
rect 15306 13550 15414 13626
rect 15786 13550 15894 13626
rect 16554 13550 16662 13626
rect 17034 13550 17142 13626
rect 17802 13550 17910 13626
rect 18282 13550 18390 13626
rect 19050 13550 19158 13626
rect 19530 13550 19638 13626
rect 20298 13550 20406 13626
rect 20778 13550 20886 13626
rect 0 13454 28 13502
rect 0 13358 28 13406
rect 330 13234 438 13310
rect 810 13234 918 13310
rect 1578 13234 1686 13310
rect 2058 13234 2166 13310
rect 2826 13234 2934 13310
rect 3306 13234 3414 13310
rect 4074 13234 4182 13310
rect 4554 13234 4662 13310
rect 5322 13234 5430 13310
rect 5802 13234 5910 13310
rect 6570 13234 6678 13310
rect 7050 13234 7158 13310
rect 7818 13234 7926 13310
rect 8298 13234 8406 13310
rect 9066 13234 9174 13310
rect 9546 13234 9654 13310
rect 10314 13234 10422 13310
rect 10794 13234 10902 13310
rect 11562 13234 11670 13310
rect 12042 13234 12150 13310
rect 12810 13234 12918 13310
rect 13290 13234 13398 13310
rect 14058 13234 14166 13310
rect 14538 13234 14646 13310
rect 15306 13234 15414 13310
rect 15786 13234 15894 13310
rect 16554 13234 16662 13310
rect 17034 13234 17142 13310
rect 17802 13234 17910 13310
rect 18282 13234 18390 13310
rect 19050 13234 19158 13310
rect 19530 13234 19638 13310
rect 20298 13234 20406 13310
rect 20778 13234 20886 13310
rect 0 13138 28 13186
rect 330 12980 438 13090
rect 810 12980 918 13090
rect 1578 12980 1686 13090
rect 2058 12980 2166 13090
rect 2826 12980 2934 13090
rect 3306 12980 3414 13090
rect 4074 12980 4182 13090
rect 4554 12980 4662 13090
rect 5322 12980 5430 13090
rect 5802 12980 5910 13090
rect 6570 12980 6678 13090
rect 7050 12980 7158 13090
rect 7818 12980 7926 13090
rect 8298 12980 8406 13090
rect 9066 12980 9174 13090
rect 9546 12980 9654 13090
rect 10314 12980 10422 13090
rect 10794 12980 10902 13090
rect 11562 12980 11670 13090
rect 12042 12980 12150 13090
rect 12810 12980 12918 13090
rect 13290 12980 13398 13090
rect 14058 12980 14166 13090
rect 14538 12980 14646 13090
rect 15306 12980 15414 13090
rect 15786 12980 15894 13090
rect 16554 12980 16662 13090
rect 17034 12980 17142 13090
rect 17802 12980 17910 13090
rect 18282 12980 18390 13090
rect 19050 12980 19158 13090
rect 19530 12980 19638 13090
rect 20298 12980 20406 13090
rect 20778 12980 20886 13090
rect 0 12884 28 12932
rect 330 12760 438 12836
rect 810 12760 918 12836
rect 1578 12760 1686 12836
rect 2058 12760 2166 12836
rect 2826 12760 2934 12836
rect 3306 12760 3414 12836
rect 4074 12760 4182 12836
rect 4554 12760 4662 12836
rect 5322 12760 5430 12836
rect 5802 12760 5910 12836
rect 6570 12760 6678 12836
rect 7050 12760 7158 12836
rect 7818 12760 7926 12836
rect 8298 12760 8406 12836
rect 9066 12760 9174 12836
rect 9546 12760 9654 12836
rect 10314 12760 10422 12836
rect 10794 12760 10902 12836
rect 11562 12760 11670 12836
rect 12042 12760 12150 12836
rect 12810 12760 12918 12836
rect 13290 12760 13398 12836
rect 14058 12760 14166 12836
rect 14538 12760 14646 12836
rect 15306 12760 15414 12836
rect 15786 12760 15894 12836
rect 16554 12760 16662 12836
rect 17034 12760 17142 12836
rect 17802 12760 17910 12836
rect 18282 12760 18390 12836
rect 19050 12760 19158 12836
rect 19530 12760 19638 12836
rect 20298 12760 20406 12836
rect 20778 12760 20886 12836
rect 0 12664 28 12712
rect 0 12568 28 12616
rect 330 12444 438 12520
rect 810 12444 918 12520
rect 1578 12444 1686 12520
rect 2058 12444 2166 12520
rect 2826 12444 2934 12520
rect 3306 12444 3414 12520
rect 4074 12444 4182 12520
rect 4554 12444 4662 12520
rect 5322 12444 5430 12520
rect 5802 12444 5910 12520
rect 6570 12444 6678 12520
rect 7050 12444 7158 12520
rect 7818 12444 7926 12520
rect 8298 12444 8406 12520
rect 9066 12444 9174 12520
rect 9546 12444 9654 12520
rect 10314 12444 10422 12520
rect 10794 12444 10902 12520
rect 11562 12444 11670 12520
rect 12042 12444 12150 12520
rect 12810 12444 12918 12520
rect 13290 12444 13398 12520
rect 14058 12444 14166 12520
rect 14538 12444 14646 12520
rect 15306 12444 15414 12520
rect 15786 12444 15894 12520
rect 16554 12444 16662 12520
rect 17034 12444 17142 12520
rect 17802 12444 17910 12520
rect 18282 12444 18390 12520
rect 19050 12444 19158 12520
rect 19530 12444 19638 12520
rect 20298 12444 20406 12520
rect 20778 12444 20886 12520
rect 0 12348 28 12396
rect 330 12190 438 12300
rect 810 12190 918 12300
rect 1578 12190 1686 12300
rect 2058 12190 2166 12300
rect 2826 12190 2934 12300
rect 3306 12190 3414 12300
rect 4074 12190 4182 12300
rect 4554 12190 4662 12300
rect 5322 12190 5430 12300
rect 5802 12190 5910 12300
rect 6570 12190 6678 12300
rect 7050 12190 7158 12300
rect 7818 12190 7926 12300
rect 8298 12190 8406 12300
rect 9066 12190 9174 12300
rect 9546 12190 9654 12300
rect 10314 12190 10422 12300
rect 10794 12190 10902 12300
rect 11562 12190 11670 12300
rect 12042 12190 12150 12300
rect 12810 12190 12918 12300
rect 13290 12190 13398 12300
rect 14058 12190 14166 12300
rect 14538 12190 14646 12300
rect 15306 12190 15414 12300
rect 15786 12190 15894 12300
rect 16554 12190 16662 12300
rect 17034 12190 17142 12300
rect 17802 12190 17910 12300
rect 18282 12190 18390 12300
rect 19050 12190 19158 12300
rect 19530 12190 19638 12300
rect 20298 12190 20406 12300
rect 20778 12190 20886 12300
rect 0 12094 28 12142
rect 330 11970 438 12046
rect 810 11970 918 12046
rect 1578 11970 1686 12046
rect 2058 11970 2166 12046
rect 2826 11970 2934 12046
rect 3306 11970 3414 12046
rect 4074 11970 4182 12046
rect 4554 11970 4662 12046
rect 5322 11970 5430 12046
rect 5802 11970 5910 12046
rect 6570 11970 6678 12046
rect 7050 11970 7158 12046
rect 7818 11970 7926 12046
rect 8298 11970 8406 12046
rect 9066 11970 9174 12046
rect 9546 11970 9654 12046
rect 10314 11970 10422 12046
rect 10794 11970 10902 12046
rect 11562 11970 11670 12046
rect 12042 11970 12150 12046
rect 12810 11970 12918 12046
rect 13290 11970 13398 12046
rect 14058 11970 14166 12046
rect 14538 11970 14646 12046
rect 15306 11970 15414 12046
rect 15786 11970 15894 12046
rect 16554 11970 16662 12046
rect 17034 11970 17142 12046
rect 17802 11970 17910 12046
rect 18282 11970 18390 12046
rect 19050 11970 19158 12046
rect 19530 11970 19638 12046
rect 20298 11970 20406 12046
rect 20778 11970 20886 12046
rect 0 11874 28 11922
rect 0 11778 28 11826
rect 330 11654 438 11730
rect 810 11654 918 11730
rect 1578 11654 1686 11730
rect 2058 11654 2166 11730
rect 2826 11654 2934 11730
rect 3306 11654 3414 11730
rect 4074 11654 4182 11730
rect 4554 11654 4662 11730
rect 5322 11654 5430 11730
rect 5802 11654 5910 11730
rect 6570 11654 6678 11730
rect 7050 11654 7158 11730
rect 7818 11654 7926 11730
rect 8298 11654 8406 11730
rect 9066 11654 9174 11730
rect 9546 11654 9654 11730
rect 10314 11654 10422 11730
rect 10794 11654 10902 11730
rect 11562 11654 11670 11730
rect 12042 11654 12150 11730
rect 12810 11654 12918 11730
rect 13290 11654 13398 11730
rect 14058 11654 14166 11730
rect 14538 11654 14646 11730
rect 15306 11654 15414 11730
rect 15786 11654 15894 11730
rect 16554 11654 16662 11730
rect 17034 11654 17142 11730
rect 17802 11654 17910 11730
rect 18282 11654 18390 11730
rect 19050 11654 19158 11730
rect 19530 11654 19638 11730
rect 20298 11654 20406 11730
rect 20778 11654 20886 11730
rect 0 11558 28 11606
rect 330 11400 438 11510
rect 810 11400 918 11510
rect 1578 11400 1686 11510
rect 2058 11400 2166 11510
rect 2826 11400 2934 11510
rect 3306 11400 3414 11510
rect 4074 11400 4182 11510
rect 4554 11400 4662 11510
rect 5322 11400 5430 11510
rect 5802 11400 5910 11510
rect 6570 11400 6678 11510
rect 7050 11400 7158 11510
rect 7818 11400 7926 11510
rect 8298 11400 8406 11510
rect 9066 11400 9174 11510
rect 9546 11400 9654 11510
rect 10314 11400 10422 11510
rect 10794 11400 10902 11510
rect 11562 11400 11670 11510
rect 12042 11400 12150 11510
rect 12810 11400 12918 11510
rect 13290 11400 13398 11510
rect 14058 11400 14166 11510
rect 14538 11400 14646 11510
rect 15306 11400 15414 11510
rect 15786 11400 15894 11510
rect 16554 11400 16662 11510
rect 17034 11400 17142 11510
rect 17802 11400 17910 11510
rect 18282 11400 18390 11510
rect 19050 11400 19158 11510
rect 19530 11400 19638 11510
rect 20298 11400 20406 11510
rect 20778 11400 20886 11510
rect 0 11304 28 11352
rect 330 11180 438 11256
rect 810 11180 918 11256
rect 1578 11180 1686 11256
rect 2058 11180 2166 11256
rect 2826 11180 2934 11256
rect 3306 11180 3414 11256
rect 4074 11180 4182 11256
rect 4554 11180 4662 11256
rect 5322 11180 5430 11256
rect 5802 11180 5910 11256
rect 6570 11180 6678 11256
rect 7050 11180 7158 11256
rect 7818 11180 7926 11256
rect 8298 11180 8406 11256
rect 9066 11180 9174 11256
rect 9546 11180 9654 11256
rect 10314 11180 10422 11256
rect 10794 11180 10902 11256
rect 11562 11180 11670 11256
rect 12042 11180 12150 11256
rect 12810 11180 12918 11256
rect 13290 11180 13398 11256
rect 14058 11180 14166 11256
rect 14538 11180 14646 11256
rect 15306 11180 15414 11256
rect 15786 11180 15894 11256
rect 16554 11180 16662 11256
rect 17034 11180 17142 11256
rect 17802 11180 17910 11256
rect 18282 11180 18390 11256
rect 19050 11180 19158 11256
rect 19530 11180 19638 11256
rect 20298 11180 20406 11256
rect 20778 11180 20886 11256
rect 0 11084 28 11132
rect 0 10988 28 11036
rect 330 10864 438 10940
rect 810 10864 918 10940
rect 1578 10864 1686 10940
rect 2058 10864 2166 10940
rect 2826 10864 2934 10940
rect 3306 10864 3414 10940
rect 4074 10864 4182 10940
rect 4554 10864 4662 10940
rect 5322 10864 5430 10940
rect 5802 10864 5910 10940
rect 6570 10864 6678 10940
rect 7050 10864 7158 10940
rect 7818 10864 7926 10940
rect 8298 10864 8406 10940
rect 9066 10864 9174 10940
rect 9546 10864 9654 10940
rect 10314 10864 10422 10940
rect 10794 10864 10902 10940
rect 11562 10864 11670 10940
rect 12042 10864 12150 10940
rect 12810 10864 12918 10940
rect 13290 10864 13398 10940
rect 14058 10864 14166 10940
rect 14538 10864 14646 10940
rect 15306 10864 15414 10940
rect 15786 10864 15894 10940
rect 16554 10864 16662 10940
rect 17034 10864 17142 10940
rect 17802 10864 17910 10940
rect 18282 10864 18390 10940
rect 19050 10864 19158 10940
rect 19530 10864 19638 10940
rect 20298 10864 20406 10940
rect 20778 10864 20886 10940
rect 0 10768 28 10816
rect 330 10610 438 10720
rect 810 10610 918 10720
rect 1578 10610 1686 10720
rect 2058 10610 2166 10720
rect 2826 10610 2934 10720
rect 3306 10610 3414 10720
rect 4074 10610 4182 10720
rect 4554 10610 4662 10720
rect 5322 10610 5430 10720
rect 5802 10610 5910 10720
rect 6570 10610 6678 10720
rect 7050 10610 7158 10720
rect 7818 10610 7926 10720
rect 8298 10610 8406 10720
rect 9066 10610 9174 10720
rect 9546 10610 9654 10720
rect 10314 10610 10422 10720
rect 10794 10610 10902 10720
rect 11562 10610 11670 10720
rect 12042 10610 12150 10720
rect 12810 10610 12918 10720
rect 13290 10610 13398 10720
rect 14058 10610 14166 10720
rect 14538 10610 14646 10720
rect 15306 10610 15414 10720
rect 15786 10610 15894 10720
rect 16554 10610 16662 10720
rect 17034 10610 17142 10720
rect 17802 10610 17910 10720
rect 18282 10610 18390 10720
rect 19050 10610 19158 10720
rect 19530 10610 19638 10720
rect 20298 10610 20406 10720
rect 20778 10610 20886 10720
rect 0 10514 28 10562
rect 330 10390 438 10466
rect 810 10390 918 10466
rect 1578 10390 1686 10466
rect 2058 10390 2166 10466
rect 2826 10390 2934 10466
rect 3306 10390 3414 10466
rect 4074 10390 4182 10466
rect 4554 10390 4662 10466
rect 5322 10390 5430 10466
rect 5802 10390 5910 10466
rect 6570 10390 6678 10466
rect 7050 10390 7158 10466
rect 7818 10390 7926 10466
rect 8298 10390 8406 10466
rect 9066 10390 9174 10466
rect 9546 10390 9654 10466
rect 10314 10390 10422 10466
rect 10794 10390 10902 10466
rect 11562 10390 11670 10466
rect 12042 10390 12150 10466
rect 12810 10390 12918 10466
rect 13290 10390 13398 10466
rect 14058 10390 14166 10466
rect 14538 10390 14646 10466
rect 15306 10390 15414 10466
rect 15786 10390 15894 10466
rect 16554 10390 16662 10466
rect 17034 10390 17142 10466
rect 17802 10390 17910 10466
rect 18282 10390 18390 10466
rect 19050 10390 19158 10466
rect 19530 10390 19638 10466
rect 20298 10390 20406 10466
rect 20778 10390 20886 10466
rect 0 10294 28 10342
rect 0 10198 28 10246
rect 330 10074 438 10150
rect 810 10074 918 10150
rect 1578 10074 1686 10150
rect 2058 10074 2166 10150
rect 2826 10074 2934 10150
rect 3306 10074 3414 10150
rect 4074 10074 4182 10150
rect 4554 10074 4662 10150
rect 5322 10074 5430 10150
rect 5802 10074 5910 10150
rect 6570 10074 6678 10150
rect 7050 10074 7158 10150
rect 7818 10074 7926 10150
rect 8298 10074 8406 10150
rect 9066 10074 9174 10150
rect 9546 10074 9654 10150
rect 10314 10074 10422 10150
rect 10794 10074 10902 10150
rect 11562 10074 11670 10150
rect 12042 10074 12150 10150
rect 12810 10074 12918 10150
rect 13290 10074 13398 10150
rect 14058 10074 14166 10150
rect 14538 10074 14646 10150
rect 15306 10074 15414 10150
rect 15786 10074 15894 10150
rect 16554 10074 16662 10150
rect 17034 10074 17142 10150
rect 17802 10074 17910 10150
rect 18282 10074 18390 10150
rect 19050 10074 19158 10150
rect 19530 10074 19638 10150
rect 20298 10074 20406 10150
rect 20778 10074 20886 10150
rect 0 9978 28 10026
rect 330 9820 438 9930
rect 810 9820 918 9930
rect 1578 9820 1686 9930
rect 2058 9820 2166 9930
rect 2826 9820 2934 9930
rect 3306 9820 3414 9930
rect 4074 9820 4182 9930
rect 4554 9820 4662 9930
rect 5322 9820 5430 9930
rect 5802 9820 5910 9930
rect 6570 9820 6678 9930
rect 7050 9820 7158 9930
rect 7818 9820 7926 9930
rect 8298 9820 8406 9930
rect 9066 9820 9174 9930
rect 9546 9820 9654 9930
rect 10314 9820 10422 9930
rect 10794 9820 10902 9930
rect 11562 9820 11670 9930
rect 12042 9820 12150 9930
rect 12810 9820 12918 9930
rect 13290 9820 13398 9930
rect 14058 9820 14166 9930
rect 14538 9820 14646 9930
rect 15306 9820 15414 9930
rect 15786 9820 15894 9930
rect 16554 9820 16662 9930
rect 17034 9820 17142 9930
rect 17802 9820 17910 9930
rect 18282 9820 18390 9930
rect 19050 9820 19158 9930
rect 19530 9820 19638 9930
rect 20298 9820 20406 9930
rect 20778 9820 20886 9930
rect 0 9724 28 9772
rect 330 9600 438 9676
rect 810 9600 918 9676
rect 1578 9600 1686 9676
rect 2058 9600 2166 9676
rect 2826 9600 2934 9676
rect 3306 9600 3414 9676
rect 4074 9600 4182 9676
rect 4554 9600 4662 9676
rect 5322 9600 5430 9676
rect 5802 9600 5910 9676
rect 6570 9600 6678 9676
rect 7050 9600 7158 9676
rect 7818 9600 7926 9676
rect 8298 9600 8406 9676
rect 9066 9600 9174 9676
rect 9546 9600 9654 9676
rect 10314 9600 10422 9676
rect 10794 9600 10902 9676
rect 11562 9600 11670 9676
rect 12042 9600 12150 9676
rect 12810 9600 12918 9676
rect 13290 9600 13398 9676
rect 14058 9600 14166 9676
rect 14538 9600 14646 9676
rect 15306 9600 15414 9676
rect 15786 9600 15894 9676
rect 16554 9600 16662 9676
rect 17034 9600 17142 9676
rect 17802 9600 17910 9676
rect 18282 9600 18390 9676
rect 19050 9600 19158 9676
rect 19530 9600 19638 9676
rect 20298 9600 20406 9676
rect 20778 9600 20886 9676
rect 0 9504 28 9552
rect 0 9408 28 9456
rect 330 9284 438 9360
rect 810 9284 918 9360
rect 1578 9284 1686 9360
rect 2058 9284 2166 9360
rect 2826 9284 2934 9360
rect 3306 9284 3414 9360
rect 4074 9284 4182 9360
rect 4554 9284 4662 9360
rect 5322 9284 5430 9360
rect 5802 9284 5910 9360
rect 6570 9284 6678 9360
rect 7050 9284 7158 9360
rect 7818 9284 7926 9360
rect 8298 9284 8406 9360
rect 9066 9284 9174 9360
rect 9546 9284 9654 9360
rect 10314 9284 10422 9360
rect 10794 9284 10902 9360
rect 11562 9284 11670 9360
rect 12042 9284 12150 9360
rect 12810 9284 12918 9360
rect 13290 9284 13398 9360
rect 14058 9284 14166 9360
rect 14538 9284 14646 9360
rect 15306 9284 15414 9360
rect 15786 9284 15894 9360
rect 16554 9284 16662 9360
rect 17034 9284 17142 9360
rect 17802 9284 17910 9360
rect 18282 9284 18390 9360
rect 19050 9284 19158 9360
rect 19530 9284 19638 9360
rect 20298 9284 20406 9360
rect 20778 9284 20886 9360
rect 0 9188 28 9236
rect 330 9030 438 9140
rect 810 9030 918 9140
rect 1578 9030 1686 9140
rect 2058 9030 2166 9140
rect 2826 9030 2934 9140
rect 3306 9030 3414 9140
rect 4074 9030 4182 9140
rect 4554 9030 4662 9140
rect 5322 9030 5430 9140
rect 5802 9030 5910 9140
rect 6570 9030 6678 9140
rect 7050 9030 7158 9140
rect 7818 9030 7926 9140
rect 8298 9030 8406 9140
rect 9066 9030 9174 9140
rect 9546 9030 9654 9140
rect 10314 9030 10422 9140
rect 10794 9030 10902 9140
rect 11562 9030 11670 9140
rect 12042 9030 12150 9140
rect 12810 9030 12918 9140
rect 13290 9030 13398 9140
rect 14058 9030 14166 9140
rect 14538 9030 14646 9140
rect 15306 9030 15414 9140
rect 15786 9030 15894 9140
rect 16554 9030 16662 9140
rect 17034 9030 17142 9140
rect 17802 9030 17910 9140
rect 18282 9030 18390 9140
rect 19050 9030 19158 9140
rect 19530 9030 19638 9140
rect 20298 9030 20406 9140
rect 20778 9030 20886 9140
rect 0 8934 28 8982
rect 330 8810 438 8886
rect 810 8810 918 8886
rect 1578 8810 1686 8886
rect 2058 8810 2166 8886
rect 2826 8810 2934 8886
rect 3306 8810 3414 8886
rect 4074 8810 4182 8886
rect 4554 8810 4662 8886
rect 5322 8810 5430 8886
rect 5802 8810 5910 8886
rect 6570 8810 6678 8886
rect 7050 8810 7158 8886
rect 7818 8810 7926 8886
rect 8298 8810 8406 8886
rect 9066 8810 9174 8886
rect 9546 8810 9654 8886
rect 10314 8810 10422 8886
rect 10794 8810 10902 8886
rect 11562 8810 11670 8886
rect 12042 8810 12150 8886
rect 12810 8810 12918 8886
rect 13290 8810 13398 8886
rect 14058 8810 14166 8886
rect 14538 8810 14646 8886
rect 15306 8810 15414 8886
rect 15786 8810 15894 8886
rect 16554 8810 16662 8886
rect 17034 8810 17142 8886
rect 17802 8810 17910 8886
rect 18282 8810 18390 8886
rect 19050 8810 19158 8886
rect 19530 8810 19638 8886
rect 20298 8810 20406 8886
rect 20778 8810 20886 8886
rect 0 8714 28 8762
rect 0 8618 28 8666
rect 330 8494 438 8570
rect 810 8494 918 8570
rect 1578 8494 1686 8570
rect 2058 8494 2166 8570
rect 2826 8494 2934 8570
rect 3306 8494 3414 8570
rect 4074 8494 4182 8570
rect 4554 8494 4662 8570
rect 5322 8494 5430 8570
rect 5802 8494 5910 8570
rect 6570 8494 6678 8570
rect 7050 8494 7158 8570
rect 7818 8494 7926 8570
rect 8298 8494 8406 8570
rect 9066 8494 9174 8570
rect 9546 8494 9654 8570
rect 10314 8494 10422 8570
rect 10794 8494 10902 8570
rect 11562 8494 11670 8570
rect 12042 8494 12150 8570
rect 12810 8494 12918 8570
rect 13290 8494 13398 8570
rect 14058 8494 14166 8570
rect 14538 8494 14646 8570
rect 15306 8494 15414 8570
rect 15786 8494 15894 8570
rect 16554 8494 16662 8570
rect 17034 8494 17142 8570
rect 17802 8494 17910 8570
rect 18282 8494 18390 8570
rect 19050 8494 19158 8570
rect 19530 8494 19638 8570
rect 20298 8494 20406 8570
rect 20778 8494 20886 8570
rect 0 8398 28 8446
rect 330 8240 438 8350
rect 810 8240 918 8350
rect 1578 8240 1686 8350
rect 2058 8240 2166 8350
rect 2826 8240 2934 8350
rect 3306 8240 3414 8350
rect 4074 8240 4182 8350
rect 4554 8240 4662 8350
rect 5322 8240 5430 8350
rect 5802 8240 5910 8350
rect 6570 8240 6678 8350
rect 7050 8240 7158 8350
rect 7818 8240 7926 8350
rect 8298 8240 8406 8350
rect 9066 8240 9174 8350
rect 9546 8240 9654 8350
rect 10314 8240 10422 8350
rect 10794 8240 10902 8350
rect 11562 8240 11670 8350
rect 12042 8240 12150 8350
rect 12810 8240 12918 8350
rect 13290 8240 13398 8350
rect 14058 8240 14166 8350
rect 14538 8240 14646 8350
rect 15306 8240 15414 8350
rect 15786 8240 15894 8350
rect 16554 8240 16662 8350
rect 17034 8240 17142 8350
rect 17802 8240 17910 8350
rect 18282 8240 18390 8350
rect 19050 8240 19158 8350
rect 19530 8240 19638 8350
rect 20298 8240 20406 8350
rect 20778 8240 20886 8350
rect 0 8144 28 8192
rect 330 8020 438 8096
rect 810 8020 918 8096
rect 1578 8020 1686 8096
rect 2058 8020 2166 8096
rect 2826 8020 2934 8096
rect 3306 8020 3414 8096
rect 4074 8020 4182 8096
rect 4554 8020 4662 8096
rect 5322 8020 5430 8096
rect 5802 8020 5910 8096
rect 6570 8020 6678 8096
rect 7050 8020 7158 8096
rect 7818 8020 7926 8096
rect 8298 8020 8406 8096
rect 9066 8020 9174 8096
rect 9546 8020 9654 8096
rect 10314 8020 10422 8096
rect 10794 8020 10902 8096
rect 11562 8020 11670 8096
rect 12042 8020 12150 8096
rect 12810 8020 12918 8096
rect 13290 8020 13398 8096
rect 14058 8020 14166 8096
rect 14538 8020 14646 8096
rect 15306 8020 15414 8096
rect 15786 8020 15894 8096
rect 16554 8020 16662 8096
rect 17034 8020 17142 8096
rect 17802 8020 17910 8096
rect 18282 8020 18390 8096
rect 19050 8020 19158 8096
rect 19530 8020 19638 8096
rect 20298 8020 20406 8096
rect 20778 8020 20886 8096
rect 0 7924 28 7972
rect 0 7828 28 7876
rect 330 7704 438 7780
rect 810 7704 918 7780
rect 1578 7704 1686 7780
rect 2058 7704 2166 7780
rect 2826 7704 2934 7780
rect 3306 7704 3414 7780
rect 4074 7704 4182 7780
rect 4554 7704 4662 7780
rect 5322 7704 5430 7780
rect 5802 7704 5910 7780
rect 6570 7704 6678 7780
rect 7050 7704 7158 7780
rect 7818 7704 7926 7780
rect 8298 7704 8406 7780
rect 9066 7704 9174 7780
rect 9546 7704 9654 7780
rect 10314 7704 10422 7780
rect 10794 7704 10902 7780
rect 11562 7704 11670 7780
rect 12042 7704 12150 7780
rect 12810 7704 12918 7780
rect 13290 7704 13398 7780
rect 14058 7704 14166 7780
rect 14538 7704 14646 7780
rect 15306 7704 15414 7780
rect 15786 7704 15894 7780
rect 16554 7704 16662 7780
rect 17034 7704 17142 7780
rect 17802 7704 17910 7780
rect 18282 7704 18390 7780
rect 19050 7704 19158 7780
rect 19530 7704 19638 7780
rect 20298 7704 20406 7780
rect 20778 7704 20886 7780
rect 0 7608 28 7656
rect 330 7450 438 7560
rect 810 7450 918 7560
rect 1578 7450 1686 7560
rect 2058 7450 2166 7560
rect 2826 7450 2934 7560
rect 3306 7450 3414 7560
rect 4074 7450 4182 7560
rect 4554 7450 4662 7560
rect 5322 7450 5430 7560
rect 5802 7450 5910 7560
rect 6570 7450 6678 7560
rect 7050 7450 7158 7560
rect 7818 7450 7926 7560
rect 8298 7450 8406 7560
rect 9066 7450 9174 7560
rect 9546 7450 9654 7560
rect 10314 7450 10422 7560
rect 10794 7450 10902 7560
rect 11562 7450 11670 7560
rect 12042 7450 12150 7560
rect 12810 7450 12918 7560
rect 13290 7450 13398 7560
rect 14058 7450 14166 7560
rect 14538 7450 14646 7560
rect 15306 7450 15414 7560
rect 15786 7450 15894 7560
rect 16554 7450 16662 7560
rect 17034 7450 17142 7560
rect 17802 7450 17910 7560
rect 18282 7450 18390 7560
rect 19050 7450 19158 7560
rect 19530 7450 19638 7560
rect 20298 7450 20406 7560
rect 20778 7450 20886 7560
rect 0 7354 28 7402
rect 330 7230 438 7306
rect 810 7230 918 7306
rect 1578 7230 1686 7306
rect 2058 7230 2166 7306
rect 2826 7230 2934 7306
rect 3306 7230 3414 7306
rect 4074 7230 4182 7306
rect 4554 7230 4662 7306
rect 5322 7230 5430 7306
rect 5802 7230 5910 7306
rect 6570 7230 6678 7306
rect 7050 7230 7158 7306
rect 7818 7230 7926 7306
rect 8298 7230 8406 7306
rect 9066 7230 9174 7306
rect 9546 7230 9654 7306
rect 10314 7230 10422 7306
rect 10794 7230 10902 7306
rect 11562 7230 11670 7306
rect 12042 7230 12150 7306
rect 12810 7230 12918 7306
rect 13290 7230 13398 7306
rect 14058 7230 14166 7306
rect 14538 7230 14646 7306
rect 15306 7230 15414 7306
rect 15786 7230 15894 7306
rect 16554 7230 16662 7306
rect 17034 7230 17142 7306
rect 17802 7230 17910 7306
rect 18282 7230 18390 7306
rect 19050 7230 19158 7306
rect 19530 7230 19638 7306
rect 20298 7230 20406 7306
rect 20778 7230 20886 7306
rect 0 7134 28 7182
rect 0 7038 28 7086
rect 330 6914 438 6990
rect 810 6914 918 6990
rect 1578 6914 1686 6990
rect 2058 6914 2166 6990
rect 2826 6914 2934 6990
rect 3306 6914 3414 6990
rect 4074 6914 4182 6990
rect 4554 6914 4662 6990
rect 5322 6914 5430 6990
rect 5802 6914 5910 6990
rect 6570 6914 6678 6990
rect 7050 6914 7158 6990
rect 7818 6914 7926 6990
rect 8298 6914 8406 6990
rect 9066 6914 9174 6990
rect 9546 6914 9654 6990
rect 10314 6914 10422 6990
rect 10794 6914 10902 6990
rect 11562 6914 11670 6990
rect 12042 6914 12150 6990
rect 12810 6914 12918 6990
rect 13290 6914 13398 6990
rect 14058 6914 14166 6990
rect 14538 6914 14646 6990
rect 15306 6914 15414 6990
rect 15786 6914 15894 6990
rect 16554 6914 16662 6990
rect 17034 6914 17142 6990
rect 17802 6914 17910 6990
rect 18282 6914 18390 6990
rect 19050 6914 19158 6990
rect 19530 6914 19638 6990
rect 20298 6914 20406 6990
rect 20778 6914 20886 6990
rect 0 6818 28 6866
rect 330 6660 438 6770
rect 810 6660 918 6770
rect 1578 6660 1686 6770
rect 2058 6660 2166 6770
rect 2826 6660 2934 6770
rect 3306 6660 3414 6770
rect 4074 6660 4182 6770
rect 4554 6660 4662 6770
rect 5322 6660 5430 6770
rect 5802 6660 5910 6770
rect 6570 6660 6678 6770
rect 7050 6660 7158 6770
rect 7818 6660 7926 6770
rect 8298 6660 8406 6770
rect 9066 6660 9174 6770
rect 9546 6660 9654 6770
rect 10314 6660 10422 6770
rect 10794 6660 10902 6770
rect 11562 6660 11670 6770
rect 12042 6660 12150 6770
rect 12810 6660 12918 6770
rect 13290 6660 13398 6770
rect 14058 6660 14166 6770
rect 14538 6660 14646 6770
rect 15306 6660 15414 6770
rect 15786 6660 15894 6770
rect 16554 6660 16662 6770
rect 17034 6660 17142 6770
rect 17802 6660 17910 6770
rect 18282 6660 18390 6770
rect 19050 6660 19158 6770
rect 19530 6660 19638 6770
rect 20298 6660 20406 6770
rect 20778 6660 20886 6770
rect 0 6564 28 6612
rect 330 6440 438 6516
rect 810 6440 918 6516
rect 1578 6440 1686 6516
rect 2058 6440 2166 6516
rect 2826 6440 2934 6516
rect 3306 6440 3414 6516
rect 4074 6440 4182 6516
rect 4554 6440 4662 6516
rect 5322 6440 5430 6516
rect 5802 6440 5910 6516
rect 6570 6440 6678 6516
rect 7050 6440 7158 6516
rect 7818 6440 7926 6516
rect 8298 6440 8406 6516
rect 9066 6440 9174 6516
rect 9546 6440 9654 6516
rect 10314 6440 10422 6516
rect 10794 6440 10902 6516
rect 11562 6440 11670 6516
rect 12042 6440 12150 6516
rect 12810 6440 12918 6516
rect 13290 6440 13398 6516
rect 14058 6440 14166 6516
rect 14538 6440 14646 6516
rect 15306 6440 15414 6516
rect 15786 6440 15894 6516
rect 16554 6440 16662 6516
rect 17034 6440 17142 6516
rect 17802 6440 17910 6516
rect 18282 6440 18390 6516
rect 19050 6440 19158 6516
rect 19530 6440 19638 6516
rect 20298 6440 20406 6516
rect 20778 6440 20886 6516
rect 0 6344 28 6392
rect 0 6248 28 6296
rect 330 6124 438 6200
rect 810 6124 918 6200
rect 1578 6124 1686 6200
rect 2058 6124 2166 6200
rect 2826 6124 2934 6200
rect 3306 6124 3414 6200
rect 4074 6124 4182 6200
rect 4554 6124 4662 6200
rect 5322 6124 5430 6200
rect 5802 6124 5910 6200
rect 6570 6124 6678 6200
rect 7050 6124 7158 6200
rect 7818 6124 7926 6200
rect 8298 6124 8406 6200
rect 9066 6124 9174 6200
rect 9546 6124 9654 6200
rect 10314 6124 10422 6200
rect 10794 6124 10902 6200
rect 11562 6124 11670 6200
rect 12042 6124 12150 6200
rect 12810 6124 12918 6200
rect 13290 6124 13398 6200
rect 14058 6124 14166 6200
rect 14538 6124 14646 6200
rect 15306 6124 15414 6200
rect 15786 6124 15894 6200
rect 16554 6124 16662 6200
rect 17034 6124 17142 6200
rect 17802 6124 17910 6200
rect 18282 6124 18390 6200
rect 19050 6124 19158 6200
rect 19530 6124 19638 6200
rect 20298 6124 20406 6200
rect 20778 6124 20886 6200
rect 0 6028 28 6076
rect 330 5870 438 5980
rect 810 5870 918 5980
rect 1578 5870 1686 5980
rect 2058 5870 2166 5980
rect 2826 5870 2934 5980
rect 3306 5870 3414 5980
rect 4074 5870 4182 5980
rect 4554 5870 4662 5980
rect 5322 5870 5430 5980
rect 5802 5870 5910 5980
rect 6570 5870 6678 5980
rect 7050 5870 7158 5980
rect 7818 5870 7926 5980
rect 8298 5870 8406 5980
rect 9066 5870 9174 5980
rect 9546 5870 9654 5980
rect 10314 5870 10422 5980
rect 10794 5870 10902 5980
rect 11562 5870 11670 5980
rect 12042 5870 12150 5980
rect 12810 5870 12918 5980
rect 13290 5870 13398 5980
rect 14058 5870 14166 5980
rect 14538 5870 14646 5980
rect 15306 5870 15414 5980
rect 15786 5870 15894 5980
rect 16554 5870 16662 5980
rect 17034 5870 17142 5980
rect 17802 5870 17910 5980
rect 18282 5870 18390 5980
rect 19050 5870 19158 5980
rect 19530 5870 19638 5980
rect 20298 5870 20406 5980
rect 20778 5870 20886 5980
rect 0 5774 28 5822
rect 330 5650 438 5726
rect 810 5650 918 5726
rect 1578 5650 1686 5726
rect 2058 5650 2166 5726
rect 2826 5650 2934 5726
rect 3306 5650 3414 5726
rect 4074 5650 4182 5726
rect 4554 5650 4662 5726
rect 5322 5650 5430 5726
rect 5802 5650 5910 5726
rect 6570 5650 6678 5726
rect 7050 5650 7158 5726
rect 7818 5650 7926 5726
rect 8298 5650 8406 5726
rect 9066 5650 9174 5726
rect 9546 5650 9654 5726
rect 10314 5650 10422 5726
rect 10794 5650 10902 5726
rect 11562 5650 11670 5726
rect 12042 5650 12150 5726
rect 12810 5650 12918 5726
rect 13290 5650 13398 5726
rect 14058 5650 14166 5726
rect 14538 5650 14646 5726
rect 15306 5650 15414 5726
rect 15786 5650 15894 5726
rect 16554 5650 16662 5726
rect 17034 5650 17142 5726
rect 17802 5650 17910 5726
rect 18282 5650 18390 5726
rect 19050 5650 19158 5726
rect 19530 5650 19638 5726
rect 20298 5650 20406 5726
rect 20778 5650 20886 5726
rect 0 5554 28 5602
rect 0 5458 28 5506
rect 330 5334 438 5410
rect 810 5334 918 5410
rect 1578 5334 1686 5410
rect 2058 5334 2166 5410
rect 2826 5334 2934 5410
rect 3306 5334 3414 5410
rect 4074 5334 4182 5410
rect 4554 5334 4662 5410
rect 5322 5334 5430 5410
rect 5802 5334 5910 5410
rect 6570 5334 6678 5410
rect 7050 5334 7158 5410
rect 7818 5334 7926 5410
rect 8298 5334 8406 5410
rect 9066 5334 9174 5410
rect 9546 5334 9654 5410
rect 10314 5334 10422 5410
rect 10794 5334 10902 5410
rect 11562 5334 11670 5410
rect 12042 5334 12150 5410
rect 12810 5334 12918 5410
rect 13290 5334 13398 5410
rect 14058 5334 14166 5410
rect 14538 5334 14646 5410
rect 15306 5334 15414 5410
rect 15786 5334 15894 5410
rect 16554 5334 16662 5410
rect 17034 5334 17142 5410
rect 17802 5334 17910 5410
rect 18282 5334 18390 5410
rect 19050 5334 19158 5410
rect 19530 5334 19638 5410
rect 20298 5334 20406 5410
rect 20778 5334 20886 5410
rect 0 5238 28 5286
rect 330 5080 438 5190
rect 810 5080 918 5190
rect 1578 5080 1686 5190
rect 2058 5080 2166 5190
rect 2826 5080 2934 5190
rect 3306 5080 3414 5190
rect 4074 5080 4182 5190
rect 4554 5080 4662 5190
rect 5322 5080 5430 5190
rect 5802 5080 5910 5190
rect 6570 5080 6678 5190
rect 7050 5080 7158 5190
rect 7818 5080 7926 5190
rect 8298 5080 8406 5190
rect 9066 5080 9174 5190
rect 9546 5080 9654 5190
rect 10314 5080 10422 5190
rect 10794 5080 10902 5190
rect 11562 5080 11670 5190
rect 12042 5080 12150 5190
rect 12810 5080 12918 5190
rect 13290 5080 13398 5190
rect 14058 5080 14166 5190
rect 14538 5080 14646 5190
rect 15306 5080 15414 5190
rect 15786 5080 15894 5190
rect 16554 5080 16662 5190
rect 17034 5080 17142 5190
rect 17802 5080 17910 5190
rect 18282 5080 18390 5190
rect 19050 5080 19158 5190
rect 19530 5080 19638 5190
rect 20298 5080 20406 5190
rect 20778 5080 20886 5190
rect 0 4984 28 5032
rect 330 4860 438 4936
rect 810 4860 918 4936
rect 1578 4860 1686 4936
rect 2058 4860 2166 4936
rect 2826 4860 2934 4936
rect 3306 4860 3414 4936
rect 4074 4860 4182 4936
rect 4554 4860 4662 4936
rect 5322 4860 5430 4936
rect 5802 4860 5910 4936
rect 6570 4860 6678 4936
rect 7050 4860 7158 4936
rect 7818 4860 7926 4936
rect 8298 4860 8406 4936
rect 9066 4860 9174 4936
rect 9546 4860 9654 4936
rect 10314 4860 10422 4936
rect 10794 4860 10902 4936
rect 11562 4860 11670 4936
rect 12042 4860 12150 4936
rect 12810 4860 12918 4936
rect 13290 4860 13398 4936
rect 14058 4860 14166 4936
rect 14538 4860 14646 4936
rect 15306 4860 15414 4936
rect 15786 4860 15894 4936
rect 16554 4860 16662 4936
rect 17034 4860 17142 4936
rect 17802 4860 17910 4936
rect 18282 4860 18390 4936
rect 19050 4860 19158 4936
rect 19530 4860 19638 4936
rect 20298 4860 20406 4936
rect 20778 4860 20886 4936
rect 0 4764 28 4812
rect 0 4668 28 4716
rect 330 4544 438 4620
rect 810 4544 918 4620
rect 1578 4544 1686 4620
rect 2058 4544 2166 4620
rect 2826 4544 2934 4620
rect 3306 4544 3414 4620
rect 4074 4544 4182 4620
rect 4554 4544 4662 4620
rect 5322 4544 5430 4620
rect 5802 4544 5910 4620
rect 6570 4544 6678 4620
rect 7050 4544 7158 4620
rect 7818 4544 7926 4620
rect 8298 4544 8406 4620
rect 9066 4544 9174 4620
rect 9546 4544 9654 4620
rect 10314 4544 10422 4620
rect 10794 4544 10902 4620
rect 11562 4544 11670 4620
rect 12042 4544 12150 4620
rect 12810 4544 12918 4620
rect 13290 4544 13398 4620
rect 14058 4544 14166 4620
rect 14538 4544 14646 4620
rect 15306 4544 15414 4620
rect 15786 4544 15894 4620
rect 16554 4544 16662 4620
rect 17034 4544 17142 4620
rect 17802 4544 17910 4620
rect 18282 4544 18390 4620
rect 19050 4544 19158 4620
rect 19530 4544 19638 4620
rect 20298 4544 20406 4620
rect 20778 4544 20886 4620
rect 0 4448 28 4496
rect 330 4290 438 4400
rect 810 4290 918 4400
rect 1578 4290 1686 4400
rect 2058 4290 2166 4400
rect 2826 4290 2934 4400
rect 3306 4290 3414 4400
rect 4074 4290 4182 4400
rect 4554 4290 4662 4400
rect 5322 4290 5430 4400
rect 5802 4290 5910 4400
rect 6570 4290 6678 4400
rect 7050 4290 7158 4400
rect 7818 4290 7926 4400
rect 8298 4290 8406 4400
rect 9066 4290 9174 4400
rect 9546 4290 9654 4400
rect 10314 4290 10422 4400
rect 10794 4290 10902 4400
rect 11562 4290 11670 4400
rect 12042 4290 12150 4400
rect 12810 4290 12918 4400
rect 13290 4290 13398 4400
rect 14058 4290 14166 4400
rect 14538 4290 14646 4400
rect 15306 4290 15414 4400
rect 15786 4290 15894 4400
rect 16554 4290 16662 4400
rect 17034 4290 17142 4400
rect 17802 4290 17910 4400
rect 18282 4290 18390 4400
rect 19050 4290 19158 4400
rect 19530 4290 19638 4400
rect 20298 4290 20406 4400
rect 20778 4290 20886 4400
rect 0 4194 28 4242
rect 330 4070 438 4146
rect 810 4070 918 4146
rect 1578 4070 1686 4146
rect 2058 4070 2166 4146
rect 2826 4070 2934 4146
rect 3306 4070 3414 4146
rect 4074 4070 4182 4146
rect 4554 4070 4662 4146
rect 5322 4070 5430 4146
rect 5802 4070 5910 4146
rect 6570 4070 6678 4146
rect 7050 4070 7158 4146
rect 7818 4070 7926 4146
rect 8298 4070 8406 4146
rect 9066 4070 9174 4146
rect 9546 4070 9654 4146
rect 10314 4070 10422 4146
rect 10794 4070 10902 4146
rect 11562 4070 11670 4146
rect 12042 4070 12150 4146
rect 12810 4070 12918 4146
rect 13290 4070 13398 4146
rect 14058 4070 14166 4146
rect 14538 4070 14646 4146
rect 15306 4070 15414 4146
rect 15786 4070 15894 4146
rect 16554 4070 16662 4146
rect 17034 4070 17142 4146
rect 17802 4070 17910 4146
rect 18282 4070 18390 4146
rect 19050 4070 19158 4146
rect 19530 4070 19638 4146
rect 20298 4070 20406 4146
rect 20778 4070 20886 4146
rect 0 3974 28 4022
rect 0 3878 28 3926
rect 330 3754 438 3830
rect 810 3754 918 3830
rect 1578 3754 1686 3830
rect 2058 3754 2166 3830
rect 2826 3754 2934 3830
rect 3306 3754 3414 3830
rect 4074 3754 4182 3830
rect 4554 3754 4662 3830
rect 5322 3754 5430 3830
rect 5802 3754 5910 3830
rect 6570 3754 6678 3830
rect 7050 3754 7158 3830
rect 7818 3754 7926 3830
rect 8298 3754 8406 3830
rect 9066 3754 9174 3830
rect 9546 3754 9654 3830
rect 10314 3754 10422 3830
rect 10794 3754 10902 3830
rect 11562 3754 11670 3830
rect 12042 3754 12150 3830
rect 12810 3754 12918 3830
rect 13290 3754 13398 3830
rect 14058 3754 14166 3830
rect 14538 3754 14646 3830
rect 15306 3754 15414 3830
rect 15786 3754 15894 3830
rect 16554 3754 16662 3830
rect 17034 3754 17142 3830
rect 17802 3754 17910 3830
rect 18282 3754 18390 3830
rect 19050 3754 19158 3830
rect 19530 3754 19638 3830
rect 20298 3754 20406 3830
rect 20778 3754 20886 3830
rect 0 3658 28 3706
rect 330 3500 438 3610
rect 810 3500 918 3610
rect 1578 3500 1686 3610
rect 2058 3500 2166 3610
rect 2826 3500 2934 3610
rect 3306 3500 3414 3610
rect 4074 3500 4182 3610
rect 4554 3500 4662 3610
rect 5322 3500 5430 3610
rect 5802 3500 5910 3610
rect 6570 3500 6678 3610
rect 7050 3500 7158 3610
rect 7818 3500 7926 3610
rect 8298 3500 8406 3610
rect 9066 3500 9174 3610
rect 9546 3500 9654 3610
rect 10314 3500 10422 3610
rect 10794 3500 10902 3610
rect 11562 3500 11670 3610
rect 12042 3500 12150 3610
rect 12810 3500 12918 3610
rect 13290 3500 13398 3610
rect 14058 3500 14166 3610
rect 14538 3500 14646 3610
rect 15306 3500 15414 3610
rect 15786 3500 15894 3610
rect 16554 3500 16662 3610
rect 17034 3500 17142 3610
rect 17802 3500 17910 3610
rect 18282 3500 18390 3610
rect 19050 3500 19158 3610
rect 19530 3500 19638 3610
rect 20298 3500 20406 3610
rect 20778 3500 20886 3610
rect 0 3404 28 3452
rect 330 3280 438 3356
rect 810 3280 918 3356
rect 1578 3280 1686 3356
rect 2058 3280 2166 3356
rect 2826 3280 2934 3356
rect 3306 3280 3414 3356
rect 4074 3280 4182 3356
rect 4554 3280 4662 3356
rect 5322 3280 5430 3356
rect 5802 3280 5910 3356
rect 6570 3280 6678 3356
rect 7050 3280 7158 3356
rect 7818 3280 7926 3356
rect 8298 3280 8406 3356
rect 9066 3280 9174 3356
rect 9546 3280 9654 3356
rect 10314 3280 10422 3356
rect 10794 3280 10902 3356
rect 11562 3280 11670 3356
rect 12042 3280 12150 3356
rect 12810 3280 12918 3356
rect 13290 3280 13398 3356
rect 14058 3280 14166 3356
rect 14538 3280 14646 3356
rect 15306 3280 15414 3356
rect 15786 3280 15894 3356
rect 16554 3280 16662 3356
rect 17034 3280 17142 3356
rect 17802 3280 17910 3356
rect 18282 3280 18390 3356
rect 19050 3280 19158 3356
rect 19530 3280 19638 3356
rect 20298 3280 20406 3356
rect 20778 3280 20886 3356
rect 0 3184 28 3232
rect 0 3088 28 3136
rect 330 2964 438 3040
rect 810 2964 918 3040
rect 1578 2964 1686 3040
rect 2058 2964 2166 3040
rect 2826 2964 2934 3040
rect 3306 2964 3414 3040
rect 4074 2964 4182 3040
rect 4554 2964 4662 3040
rect 5322 2964 5430 3040
rect 5802 2964 5910 3040
rect 6570 2964 6678 3040
rect 7050 2964 7158 3040
rect 7818 2964 7926 3040
rect 8298 2964 8406 3040
rect 9066 2964 9174 3040
rect 9546 2964 9654 3040
rect 10314 2964 10422 3040
rect 10794 2964 10902 3040
rect 11562 2964 11670 3040
rect 12042 2964 12150 3040
rect 12810 2964 12918 3040
rect 13290 2964 13398 3040
rect 14058 2964 14166 3040
rect 14538 2964 14646 3040
rect 15306 2964 15414 3040
rect 15786 2964 15894 3040
rect 16554 2964 16662 3040
rect 17034 2964 17142 3040
rect 17802 2964 17910 3040
rect 18282 2964 18390 3040
rect 19050 2964 19158 3040
rect 19530 2964 19638 3040
rect 20298 2964 20406 3040
rect 20778 2964 20886 3040
rect 0 2868 28 2916
rect 330 2710 438 2820
rect 810 2710 918 2820
rect 1578 2710 1686 2820
rect 2058 2710 2166 2820
rect 2826 2710 2934 2820
rect 3306 2710 3414 2820
rect 4074 2710 4182 2820
rect 4554 2710 4662 2820
rect 5322 2710 5430 2820
rect 5802 2710 5910 2820
rect 6570 2710 6678 2820
rect 7050 2710 7158 2820
rect 7818 2710 7926 2820
rect 8298 2710 8406 2820
rect 9066 2710 9174 2820
rect 9546 2710 9654 2820
rect 10314 2710 10422 2820
rect 10794 2710 10902 2820
rect 11562 2710 11670 2820
rect 12042 2710 12150 2820
rect 12810 2710 12918 2820
rect 13290 2710 13398 2820
rect 14058 2710 14166 2820
rect 14538 2710 14646 2820
rect 15306 2710 15414 2820
rect 15786 2710 15894 2820
rect 16554 2710 16662 2820
rect 17034 2710 17142 2820
rect 17802 2710 17910 2820
rect 18282 2710 18390 2820
rect 19050 2710 19158 2820
rect 19530 2710 19638 2820
rect 20298 2710 20406 2820
rect 20778 2710 20886 2820
rect 0 2614 28 2662
rect 330 2490 438 2566
rect 810 2490 918 2566
rect 1578 2490 1686 2566
rect 2058 2490 2166 2566
rect 2826 2490 2934 2566
rect 3306 2490 3414 2566
rect 4074 2490 4182 2566
rect 4554 2490 4662 2566
rect 5322 2490 5430 2566
rect 5802 2490 5910 2566
rect 6570 2490 6678 2566
rect 7050 2490 7158 2566
rect 7818 2490 7926 2566
rect 8298 2490 8406 2566
rect 9066 2490 9174 2566
rect 9546 2490 9654 2566
rect 10314 2490 10422 2566
rect 10794 2490 10902 2566
rect 11562 2490 11670 2566
rect 12042 2490 12150 2566
rect 12810 2490 12918 2566
rect 13290 2490 13398 2566
rect 14058 2490 14166 2566
rect 14538 2490 14646 2566
rect 15306 2490 15414 2566
rect 15786 2490 15894 2566
rect 16554 2490 16662 2566
rect 17034 2490 17142 2566
rect 17802 2490 17910 2566
rect 18282 2490 18390 2566
rect 19050 2490 19158 2566
rect 19530 2490 19638 2566
rect 20298 2490 20406 2566
rect 20778 2490 20886 2566
rect 0 2394 28 2442
rect 0 2298 28 2346
rect 330 2174 438 2250
rect 810 2174 918 2250
rect 1578 2174 1686 2250
rect 2058 2174 2166 2250
rect 2826 2174 2934 2250
rect 3306 2174 3414 2250
rect 4074 2174 4182 2250
rect 4554 2174 4662 2250
rect 5322 2174 5430 2250
rect 5802 2174 5910 2250
rect 6570 2174 6678 2250
rect 7050 2174 7158 2250
rect 7818 2174 7926 2250
rect 8298 2174 8406 2250
rect 9066 2174 9174 2250
rect 9546 2174 9654 2250
rect 10314 2174 10422 2250
rect 10794 2174 10902 2250
rect 11562 2174 11670 2250
rect 12042 2174 12150 2250
rect 12810 2174 12918 2250
rect 13290 2174 13398 2250
rect 14058 2174 14166 2250
rect 14538 2174 14646 2250
rect 15306 2174 15414 2250
rect 15786 2174 15894 2250
rect 16554 2174 16662 2250
rect 17034 2174 17142 2250
rect 17802 2174 17910 2250
rect 18282 2174 18390 2250
rect 19050 2174 19158 2250
rect 19530 2174 19638 2250
rect 20298 2174 20406 2250
rect 20778 2174 20886 2250
rect 0 2078 28 2126
rect 330 1920 438 2030
rect 810 1920 918 2030
rect 1578 1920 1686 2030
rect 2058 1920 2166 2030
rect 2826 1920 2934 2030
rect 3306 1920 3414 2030
rect 4074 1920 4182 2030
rect 4554 1920 4662 2030
rect 5322 1920 5430 2030
rect 5802 1920 5910 2030
rect 6570 1920 6678 2030
rect 7050 1920 7158 2030
rect 7818 1920 7926 2030
rect 8298 1920 8406 2030
rect 9066 1920 9174 2030
rect 9546 1920 9654 2030
rect 10314 1920 10422 2030
rect 10794 1920 10902 2030
rect 11562 1920 11670 2030
rect 12042 1920 12150 2030
rect 12810 1920 12918 2030
rect 13290 1920 13398 2030
rect 14058 1920 14166 2030
rect 14538 1920 14646 2030
rect 15306 1920 15414 2030
rect 15786 1920 15894 2030
rect 16554 1920 16662 2030
rect 17034 1920 17142 2030
rect 17802 1920 17910 2030
rect 18282 1920 18390 2030
rect 19050 1920 19158 2030
rect 19530 1920 19638 2030
rect 20298 1920 20406 2030
rect 20778 1920 20886 2030
rect 0 1824 28 1872
rect 330 1700 438 1776
rect 810 1700 918 1776
rect 1578 1700 1686 1776
rect 2058 1700 2166 1776
rect 2826 1700 2934 1776
rect 3306 1700 3414 1776
rect 4074 1700 4182 1776
rect 4554 1700 4662 1776
rect 5322 1700 5430 1776
rect 5802 1700 5910 1776
rect 6570 1700 6678 1776
rect 7050 1700 7158 1776
rect 7818 1700 7926 1776
rect 8298 1700 8406 1776
rect 9066 1700 9174 1776
rect 9546 1700 9654 1776
rect 10314 1700 10422 1776
rect 10794 1700 10902 1776
rect 11562 1700 11670 1776
rect 12042 1700 12150 1776
rect 12810 1700 12918 1776
rect 13290 1700 13398 1776
rect 14058 1700 14166 1776
rect 14538 1700 14646 1776
rect 15306 1700 15414 1776
rect 15786 1700 15894 1776
rect 16554 1700 16662 1776
rect 17034 1700 17142 1776
rect 17802 1700 17910 1776
rect 18282 1700 18390 1776
rect 19050 1700 19158 1776
rect 19530 1700 19638 1776
rect 20298 1700 20406 1776
rect 20778 1700 20886 1776
rect 0 1604 28 1652
rect 0 1508 28 1556
rect 330 1384 438 1460
rect 810 1384 918 1460
rect 1578 1384 1686 1460
rect 2058 1384 2166 1460
rect 2826 1384 2934 1460
rect 3306 1384 3414 1460
rect 4074 1384 4182 1460
rect 4554 1384 4662 1460
rect 5322 1384 5430 1460
rect 5802 1384 5910 1460
rect 6570 1384 6678 1460
rect 7050 1384 7158 1460
rect 7818 1384 7926 1460
rect 8298 1384 8406 1460
rect 9066 1384 9174 1460
rect 9546 1384 9654 1460
rect 10314 1384 10422 1460
rect 10794 1384 10902 1460
rect 11562 1384 11670 1460
rect 12042 1384 12150 1460
rect 12810 1384 12918 1460
rect 13290 1384 13398 1460
rect 14058 1384 14166 1460
rect 14538 1384 14646 1460
rect 15306 1384 15414 1460
rect 15786 1384 15894 1460
rect 16554 1384 16662 1460
rect 17034 1384 17142 1460
rect 17802 1384 17910 1460
rect 18282 1384 18390 1460
rect 19050 1384 19158 1460
rect 19530 1384 19638 1460
rect 20298 1384 20406 1460
rect 20778 1384 20886 1460
rect 0 1288 28 1336
rect 330 1130 438 1240
rect 810 1130 918 1240
rect 1578 1130 1686 1240
rect 2058 1130 2166 1240
rect 2826 1130 2934 1240
rect 3306 1130 3414 1240
rect 4074 1130 4182 1240
rect 4554 1130 4662 1240
rect 5322 1130 5430 1240
rect 5802 1130 5910 1240
rect 6570 1130 6678 1240
rect 7050 1130 7158 1240
rect 7818 1130 7926 1240
rect 8298 1130 8406 1240
rect 9066 1130 9174 1240
rect 9546 1130 9654 1240
rect 10314 1130 10422 1240
rect 10794 1130 10902 1240
rect 11562 1130 11670 1240
rect 12042 1130 12150 1240
rect 12810 1130 12918 1240
rect 13290 1130 13398 1240
rect 14058 1130 14166 1240
rect 14538 1130 14646 1240
rect 15306 1130 15414 1240
rect 15786 1130 15894 1240
rect 16554 1130 16662 1240
rect 17034 1130 17142 1240
rect 17802 1130 17910 1240
rect 18282 1130 18390 1240
rect 19050 1130 19158 1240
rect 19530 1130 19638 1240
rect 20298 1130 20406 1240
rect 20778 1130 20886 1240
rect 0 1034 28 1082
rect 330 910 438 986
rect 810 910 918 986
rect 1578 910 1686 986
rect 2058 910 2166 986
rect 2826 910 2934 986
rect 3306 910 3414 986
rect 4074 910 4182 986
rect 4554 910 4662 986
rect 5322 910 5430 986
rect 5802 910 5910 986
rect 6570 910 6678 986
rect 7050 910 7158 986
rect 7818 910 7926 986
rect 8298 910 8406 986
rect 9066 910 9174 986
rect 9546 910 9654 986
rect 10314 910 10422 986
rect 10794 910 10902 986
rect 11562 910 11670 986
rect 12042 910 12150 986
rect 12810 910 12918 986
rect 13290 910 13398 986
rect 14058 910 14166 986
rect 14538 910 14646 986
rect 15306 910 15414 986
rect 15786 910 15894 986
rect 16554 910 16662 986
rect 17034 910 17142 986
rect 17802 910 17910 986
rect 18282 910 18390 986
rect 19050 910 19158 986
rect 19530 910 19638 986
rect 20298 910 20406 986
rect 20778 910 20886 986
rect 0 814 28 862
rect 0 718 28 766
rect 330 594 438 670
rect 810 594 918 670
rect 1578 594 1686 670
rect 2058 594 2166 670
rect 2826 594 2934 670
rect 3306 594 3414 670
rect 4074 594 4182 670
rect 4554 594 4662 670
rect 5322 594 5430 670
rect 5802 594 5910 670
rect 6570 594 6678 670
rect 7050 594 7158 670
rect 7818 594 7926 670
rect 8298 594 8406 670
rect 9066 594 9174 670
rect 9546 594 9654 670
rect 10314 594 10422 670
rect 10794 594 10902 670
rect 11562 594 11670 670
rect 12042 594 12150 670
rect 12810 594 12918 670
rect 13290 594 13398 670
rect 14058 594 14166 670
rect 14538 594 14646 670
rect 15306 594 15414 670
rect 15786 594 15894 670
rect 16554 594 16662 670
rect 17034 594 17142 670
rect 17802 594 17910 670
rect 18282 594 18390 670
rect 19050 594 19158 670
rect 19530 594 19638 670
rect 20298 594 20406 670
rect 20778 594 20886 670
rect 0 498 28 546
rect 330 340 438 450
rect 810 340 918 450
rect 1578 340 1686 450
rect 2058 340 2166 450
rect 2826 340 2934 450
rect 3306 340 3414 450
rect 4074 340 4182 450
rect 4554 340 4662 450
rect 5322 340 5430 450
rect 5802 340 5910 450
rect 6570 340 6678 450
rect 7050 340 7158 450
rect 7818 340 7926 450
rect 8298 340 8406 450
rect 9066 340 9174 450
rect 9546 340 9654 450
rect 10314 340 10422 450
rect 10794 340 10902 450
rect 11562 340 11670 450
rect 12042 340 12150 450
rect 12810 340 12918 450
rect 13290 340 13398 450
rect 14058 340 14166 450
rect 14538 340 14646 450
rect 15306 340 15414 450
rect 15786 340 15894 450
rect 16554 340 16662 450
rect 17034 340 17142 450
rect 17802 340 17910 450
rect 18282 340 18390 450
rect 19050 340 19158 450
rect 19530 340 19638 450
rect 20298 340 20406 450
rect 20778 340 20886 450
rect 0 244 28 292
rect 330 120 438 196
rect 810 120 918 196
rect 1578 120 1686 196
rect 2058 120 2166 196
rect 2826 120 2934 196
rect 3306 120 3414 196
rect 4074 120 4182 196
rect 4554 120 4662 196
rect 5322 120 5430 196
rect 5802 120 5910 196
rect 6570 120 6678 196
rect 7050 120 7158 196
rect 7818 120 7926 196
rect 8298 120 8406 196
rect 9066 120 9174 196
rect 9546 120 9654 196
rect 10314 120 10422 196
rect 10794 120 10902 196
rect 11562 120 11670 196
rect 12042 120 12150 196
rect 12810 120 12918 196
rect 13290 120 13398 196
rect 14058 120 14166 196
rect 14538 120 14646 196
rect 15306 120 15414 196
rect 15786 120 15894 196
rect 16554 120 16662 196
rect 17034 120 17142 196
rect 17802 120 17910 196
rect 18282 120 18390 196
rect 19050 120 19158 196
rect 19530 120 19638 196
rect 20298 120 20406 196
rect 20778 120 20886 196
rect 0 24 28 72
use subbyte2_bitcell_array  subbyte2_bitcell_array_0
timestamp 1543373562
transform 1 0 624 0 1 395
box -42 -105 20010 25385
use subbyte2_dummy_array  subbyte2_dummy_array_0
timestamp 1543373568
transform 1 0 624 0 1 25675
box -42 -105 20010 421
use subbyte2_dummy_array  subbyte2_dummy_array_1
timestamp 1543373568
transform 1 0 624 0 -1 395
box -42 -105 20010 421
use subbyte2_replica_column  subbyte2_replica_column_0
timestamp 1543373567
transform 1 0 0 0 1 0
box -26 -26 666 26096
use subbyte2_replica_column_0  subbyte2_replica_column_0_0
timestamp 1543373568
transform 1 0 20592 0 1 0
box -42 -26 650 26096
<< labels >>
rlabel metal2 s 0 718 28 766 4 wl_0_0
port 3 nsew
rlabel metal2 s 0 498 28 546 4 wl_1_0
port 5 nsew
rlabel metal2 s 0 814 28 862 4 wl_0_1
port 7 nsew
rlabel metal2 s 0 1034 28 1082 4 wl_1_1
port 9 nsew
rlabel metal2 s 0 1508 28 1556 4 wl_0_2
port 11 nsew
rlabel metal2 s 0 1288 28 1336 4 wl_1_2
port 13 nsew
rlabel metal2 s 0 1604 28 1652 4 wl_0_3
port 15 nsew
rlabel metal2 s 0 1824 28 1872 4 wl_1_3
port 17 nsew
rlabel metal2 s 0 2298 28 2346 4 wl_0_4
port 19 nsew
rlabel metal2 s 0 2078 28 2126 4 wl_1_4
port 21 nsew
rlabel metal2 s 0 2394 28 2442 4 wl_0_5
port 23 nsew
rlabel metal2 s 0 2614 28 2662 4 wl_1_5
port 25 nsew
rlabel metal2 s 0 3088 28 3136 4 wl_0_6
port 27 nsew
rlabel metal2 s 0 2868 28 2916 4 wl_1_6
port 29 nsew
rlabel metal2 s 0 3184 28 3232 4 wl_0_7
port 31 nsew
rlabel metal2 s 0 3404 28 3452 4 wl_1_7
port 33 nsew
rlabel metal2 s 0 3878 28 3926 4 wl_0_8
port 35 nsew
rlabel metal2 s 0 3658 28 3706 4 wl_1_8
port 37 nsew
rlabel metal2 s 0 3974 28 4022 4 wl_0_9
port 39 nsew
rlabel metal2 s 0 4194 28 4242 4 wl_1_9
port 41 nsew
rlabel metal2 s 0 4668 28 4716 4 wl_0_10
port 43 nsew
rlabel metal2 s 0 4448 28 4496 4 wl_1_10
port 45 nsew
rlabel metal2 s 0 4764 28 4812 4 wl_0_11
port 47 nsew
rlabel metal2 s 0 4984 28 5032 4 wl_1_11
port 49 nsew
rlabel metal2 s 0 5458 28 5506 4 wl_0_12
port 51 nsew
rlabel metal2 s 0 5238 28 5286 4 wl_1_12
port 53 nsew
rlabel metal2 s 0 5554 28 5602 4 wl_0_13
port 55 nsew
rlabel metal2 s 0 5774 28 5822 4 wl_1_13
port 57 nsew
rlabel metal2 s 0 6248 28 6296 4 wl_0_14
port 59 nsew
rlabel metal2 s 0 6028 28 6076 4 wl_1_14
port 61 nsew
rlabel metal2 s 0 6344 28 6392 4 wl_0_15
port 63 nsew
rlabel metal2 s 0 6564 28 6612 4 wl_1_15
port 65 nsew
rlabel metal2 s 0 7038 28 7086 4 wl_0_16
port 67 nsew
rlabel metal2 s 0 6818 28 6866 4 wl_1_16
port 69 nsew
rlabel metal2 s 0 7134 28 7182 4 wl_0_17
port 71 nsew
rlabel metal2 s 0 7354 28 7402 4 wl_1_17
port 73 nsew
rlabel metal2 s 0 7828 28 7876 4 wl_0_18
port 75 nsew
rlabel metal2 s 0 7608 28 7656 4 wl_1_18
port 77 nsew
rlabel metal2 s 0 7924 28 7972 4 wl_0_19
port 79 nsew
rlabel metal2 s 0 8144 28 8192 4 wl_1_19
port 81 nsew
rlabel metal2 s 0 8618 28 8666 4 wl_0_20
port 83 nsew
rlabel metal2 s 0 8398 28 8446 4 wl_1_20
port 85 nsew
rlabel metal2 s 0 8714 28 8762 4 wl_0_21
port 87 nsew
rlabel metal2 s 0 8934 28 8982 4 wl_1_21
port 89 nsew
rlabel metal2 s 0 9408 28 9456 4 wl_0_22
port 91 nsew
rlabel metal2 s 0 9188 28 9236 4 wl_1_22
port 93 nsew
rlabel metal2 s 0 9504 28 9552 4 wl_0_23
port 95 nsew
rlabel metal2 s 0 9724 28 9772 4 wl_1_23
port 97 nsew
rlabel metal2 s 0 10198 28 10246 4 wl_0_24
port 99 nsew
rlabel metal2 s 0 9978 28 10026 4 wl_1_24
port 101 nsew
rlabel metal2 s 0 10294 28 10342 4 wl_0_25
port 103 nsew
rlabel metal2 s 0 10514 28 10562 4 wl_1_25
port 105 nsew
rlabel metal2 s 0 10988 28 11036 4 wl_0_26
port 107 nsew
rlabel metal2 s 0 10768 28 10816 4 wl_1_26
port 109 nsew
rlabel metal2 s 0 11084 28 11132 4 wl_0_27
port 111 nsew
rlabel metal2 s 0 11304 28 11352 4 wl_1_27
port 113 nsew
rlabel metal2 s 0 11778 28 11826 4 wl_0_28
port 115 nsew
rlabel metal2 s 0 11558 28 11606 4 wl_1_28
port 117 nsew
rlabel metal2 s 0 11874 28 11922 4 wl_0_29
port 119 nsew
rlabel metal2 s 0 12094 28 12142 4 wl_1_29
port 121 nsew
rlabel metal2 s 0 12568 28 12616 4 wl_0_30
port 123 nsew
rlabel metal2 s 0 12348 28 12396 4 wl_1_30
port 125 nsew
rlabel metal2 s 0 12664 28 12712 4 wl_0_31
port 127 nsew
rlabel metal2 s 0 12884 28 12932 4 wl_1_31
port 129 nsew
rlabel metal2 s 0 13358 28 13406 4 wl_0_32
port 131 nsew
rlabel metal2 s 0 13138 28 13186 4 wl_1_32
port 133 nsew
rlabel metal2 s 0 13454 28 13502 4 wl_0_33
port 135 nsew
rlabel metal2 s 0 13674 28 13722 4 wl_1_33
port 137 nsew
rlabel metal2 s 0 14148 28 14196 4 wl_0_34
port 139 nsew
rlabel metal2 s 0 13928 28 13976 4 wl_1_34
port 141 nsew
rlabel metal2 s 0 14244 28 14292 4 wl_0_35
port 143 nsew
rlabel metal2 s 0 14464 28 14512 4 wl_1_35
port 145 nsew
rlabel metal2 s 0 14938 28 14986 4 wl_0_36
port 147 nsew
rlabel metal2 s 0 14718 28 14766 4 wl_1_36
port 149 nsew
rlabel metal2 s 0 15034 28 15082 4 wl_0_37
port 151 nsew
rlabel metal2 s 0 15254 28 15302 4 wl_1_37
port 153 nsew
rlabel metal2 s 0 15728 28 15776 4 wl_0_38
port 155 nsew
rlabel metal2 s 0 15508 28 15556 4 wl_1_38
port 157 nsew
rlabel metal2 s 0 15824 28 15872 4 wl_0_39
port 159 nsew
rlabel metal2 s 0 16044 28 16092 4 wl_1_39
port 161 nsew
rlabel metal2 s 0 16518 28 16566 4 wl_0_40
port 163 nsew
rlabel metal2 s 0 16298 28 16346 4 wl_1_40
port 165 nsew
rlabel metal2 s 0 16614 28 16662 4 wl_0_41
port 167 nsew
rlabel metal2 s 0 16834 28 16882 4 wl_1_41
port 169 nsew
rlabel metal2 s 0 17308 28 17356 4 wl_0_42
port 171 nsew
rlabel metal2 s 0 17088 28 17136 4 wl_1_42
port 173 nsew
rlabel metal2 s 0 17404 28 17452 4 wl_0_43
port 175 nsew
rlabel metal2 s 0 17624 28 17672 4 wl_1_43
port 177 nsew
rlabel metal2 s 0 18098 28 18146 4 wl_0_44
port 179 nsew
rlabel metal2 s 0 17878 28 17926 4 wl_1_44
port 181 nsew
rlabel metal2 s 0 18194 28 18242 4 wl_0_45
port 183 nsew
rlabel metal2 s 0 18414 28 18462 4 wl_1_45
port 185 nsew
rlabel metal2 s 0 18888 28 18936 4 wl_0_46
port 187 nsew
rlabel metal2 s 0 18668 28 18716 4 wl_1_46
port 189 nsew
rlabel metal2 s 0 18984 28 19032 4 wl_0_47
port 191 nsew
rlabel metal2 s 0 19204 28 19252 4 wl_1_47
port 193 nsew
rlabel metal2 s 0 19678 28 19726 4 wl_0_48
port 195 nsew
rlabel metal2 s 0 19458 28 19506 4 wl_1_48
port 197 nsew
rlabel metal2 s 0 19774 28 19822 4 wl_0_49
port 199 nsew
rlabel metal2 s 0 19994 28 20042 4 wl_1_49
port 201 nsew
rlabel metal2 s 0 20468 28 20516 4 wl_0_50
port 203 nsew
rlabel metal2 s 0 20248 28 20296 4 wl_1_50
port 205 nsew
rlabel metal2 s 0 20564 28 20612 4 wl_0_51
port 207 nsew
rlabel metal2 s 0 20784 28 20832 4 wl_1_51
port 209 nsew
rlabel metal2 s 0 21258 28 21306 4 wl_0_52
port 211 nsew
rlabel metal2 s 0 21038 28 21086 4 wl_1_52
port 213 nsew
rlabel metal2 s 0 21354 28 21402 4 wl_0_53
port 215 nsew
rlabel metal2 s 0 21574 28 21622 4 wl_1_53
port 217 nsew
rlabel metal2 s 0 22048 28 22096 4 wl_0_54
port 219 nsew
rlabel metal2 s 0 21828 28 21876 4 wl_1_54
port 221 nsew
rlabel metal2 s 0 22144 28 22192 4 wl_0_55
port 223 nsew
rlabel metal2 s 0 22364 28 22412 4 wl_1_55
port 225 nsew
rlabel metal2 s 0 22838 28 22886 4 wl_0_56
port 227 nsew
rlabel metal2 s 0 22618 28 22666 4 wl_1_56
port 229 nsew
rlabel metal2 s 0 22934 28 22982 4 wl_0_57
port 231 nsew
rlabel metal2 s 0 23154 28 23202 4 wl_1_57
port 233 nsew
rlabel metal2 s 0 23628 28 23676 4 wl_0_58
port 235 nsew
rlabel metal2 s 0 23408 28 23456 4 wl_1_58
port 237 nsew
rlabel metal2 s 0 23724 28 23772 4 wl_0_59
port 239 nsew
rlabel metal2 s 0 23944 28 23992 4 wl_1_59
port 241 nsew
rlabel metal2 s 0 24418 28 24466 4 wl_0_60
port 243 nsew
rlabel metal2 s 0 24198 28 24246 4 wl_1_60
port 245 nsew
rlabel metal2 s 0 24514 28 24562 4 wl_0_61
port 247 nsew
rlabel metal2 s 0 24734 28 24782 4 wl_1_61
port 249 nsew
rlabel metal2 s 0 25208 28 25256 4 wl_0_62
port 251 nsew
rlabel metal2 s 0 24988 28 25036 4 wl_1_62
port 253 nsew
rlabel metal2 s 0 25304 28 25352 4 wl_0_63
port 255 nsew
rlabel metal2 s 0 25524 28 25572 4 wl_1_63
port 257 nsew
rlabel metal2 s 0 24 28 72 4 rbl_wl_0_0
port 259 nsew
rlabel metal2 s 0 244 28 292 4 rbl_wl_0_1
port 261 nsew
rlabel metal2 s 0 25998 28 26046 4 rbl_wl_1_0
port 263 nsew
rlabel metal2 s 0 25778 28 25826 4 rbl_wl_1_1
port 265 nsew
rlabel metal1 s 702 0 738 28 4 bl_0_0
port 267 nsew
rlabel metal1 s 918 0 954 28 4 bl_1_0
port 269 nsew
rlabel metal1 s 774 0 810 28 4 br_0_0
port 271 nsew
rlabel metal1 s 990 0 1026 28 4 br_1_0
port 273 nsew
rlabel metal1 s 1758 0 1794 28 4 bl_0_1
port 275 nsew
rlabel metal1 s 1542 0 1578 28 4 bl_1_1
port 277 nsew
rlabel metal1 s 1686 0 1722 28 4 br_0_1
port 279 nsew
rlabel metal1 s 1470 0 1506 28 4 br_1_1
port 281 nsew
rlabel metal1 s 1950 0 1986 28 4 bl_0_2
port 283 nsew
rlabel metal1 s 2166 0 2202 28 4 bl_1_2
port 285 nsew
rlabel metal1 s 2022 0 2058 28 4 br_0_2
port 287 nsew
rlabel metal1 s 2238 0 2274 28 4 br_1_2
port 289 nsew
rlabel metal1 s 3006 0 3042 28 4 bl_0_3
port 291 nsew
rlabel metal1 s 2790 0 2826 28 4 bl_1_3
port 293 nsew
rlabel metal1 s 2934 0 2970 28 4 br_0_3
port 295 nsew
rlabel metal1 s 2718 0 2754 28 4 br_1_3
port 297 nsew
rlabel metal1 s 3198 0 3234 28 4 bl_0_4
port 299 nsew
rlabel metal1 s 3414 0 3450 28 4 bl_1_4
port 301 nsew
rlabel metal1 s 3270 0 3306 28 4 br_0_4
port 303 nsew
rlabel metal1 s 3486 0 3522 28 4 br_1_4
port 305 nsew
rlabel metal1 s 4254 0 4290 28 4 bl_0_5
port 307 nsew
rlabel metal1 s 4038 0 4074 28 4 bl_1_5
port 309 nsew
rlabel metal1 s 4182 0 4218 28 4 br_0_5
port 311 nsew
rlabel metal1 s 3966 0 4002 28 4 br_1_5
port 313 nsew
rlabel metal1 s 4446 0 4482 28 4 bl_0_6
port 315 nsew
rlabel metal1 s 4662 0 4698 28 4 bl_1_6
port 317 nsew
rlabel metal1 s 4518 0 4554 28 4 br_0_6
port 319 nsew
rlabel metal1 s 4734 0 4770 28 4 br_1_6
port 321 nsew
rlabel metal1 s 5502 0 5538 28 4 bl_0_7
port 323 nsew
rlabel metal1 s 5286 0 5322 28 4 bl_1_7
port 325 nsew
rlabel metal1 s 5430 0 5466 28 4 br_0_7
port 327 nsew
rlabel metal1 s 5214 0 5250 28 4 br_1_7
port 329 nsew
rlabel metal1 s 5694 0 5730 28 4 bl_0_8
port 331 nsew
rlabel metal1 s 5910 0 5946 28 4 bl_1_8
port 333 nsew
rlabel metal1 s 5766 0 5802 28 4 br_0_8
port 335 nsew
rlabel metal1 s 5982 0 6018 28 4 br_1_8
port 337 nsew
rlabel metal1 s 6750 0 6786 28 4 bl_0_9
port 339 nsew
rlabel metal1 s 6534 0 6570 28 4 bl_1_9
port 341 nsew
rlabel metal1 s 6678 0 6714 28 4 br_0_9
port 343 nsew
rlabel metal1 s 6462 0 6498 28 4 br_1_9
port 345 nsew
rlabel metal1 s 6942 0 6978 28 4 bl_0_10
port 347 nsew
rlabel metal1 s 7158 0 7194 28 4 bl_1_10
port 349 nsew
rlabel metal1 s 7014 0 7050 28 4 br_0_10
port 351 nsew
rlabel metal1 s 7230 0 7266 28 4 br_1_10
port 353 nsew
rlabel metal1 s 7998 0 8034 28 4 bl_0_11
port 355 nsew
rlabel metal1 s 7782 0 7818 28 4 bl_1_11
port 357 nsew
rlabel metal1 s 7926 0 7962 28 4 br_0_11
port 359 nsew
rlabel metal1 s 7710 0 7746 28 4 br_1_11
port 361 nsew
rlabel metal1 s 8190 0 8226 28 4 bl_0_12
port 363 nsew
rlabel metal1 s 8406 0 8442 28 4 bl_1_12
port 365 nsew
rlabel metal1 s 8262 0 8298 28 4 br_0_12
port 367 nsew
rlabel metal1 s 8478 0 8514 28 4 br_1_12
port 369 nsew
rlabel metal1 s 9246 0 9282 28 4 bl_0_13
port 371 nsew
rlabel metal1 s 9030 0 9066 28 4 bl_1_13
port 373 nsew
rlabel metal1 s 9174 0 9210 28 4 br_0_13
port 375 nsew
rlabel metal1 s 8958 0 8994 28 4 br_1_13
port 377 nsew
rlabel metal1 s 9438 0 9474 28 4 bl_0_14
port 379 nsew
rlabel metal1 s 9654 0 9690 28 4 bl_1_14
port 381 nsew
rlabel metal1 s 9510 0 9546 28 4 br_0_14
port 383 nsew
rlabel metal1 s 9726 0 9762 28 4 br_1_14
port 385 nsew
rlabel metal1 s 10494 0 10530 28 4 bl_0_15
port 387 nsew
rlabel metal1 s 10278 0 10314 28 4 bl_1_15
port 389 nsew
rlabel metal1 s 10422 0 10458 28 4 br_0_15
port 391 nsew
rlabel metal1 s 10206 0 10242 28 4 br_1_15
port 393 nsew
rlabel metal1 s 10686 0 10722 28 4 bl_0_16
port 395 nsew
rlabel metal1 s 10902 0 10938 28 4 bl_1_16
port 397 nsew
rlabel metal1 s 10758 0 10794 28 4 br_0_16
port 399 nsew
rlabel metal1 s 10974 0 11010 28 4 br_1_16
port 401 nsew
rlabel metal1 s 11742 0 11778 28 4 bl_0_17
port 403 nsew
rlabel metal1 s 11526 0 11562 28 4 bl_1_17
port 405 nsew
rlabel metal1 s 11670 0 11706 28 4 br_0_17
port 407 nsew
rlabel metal1 s 11454 0 11490 28 4 br_1_17
port 409 nsew
rlabel metal1 s 11934 0 11970 28 4 bl_0_18
port 411 nsew
rlabel metal1 s 12150 0 12186 28 4 bl_1_18
port 413 nsew
rlabel metal1 s 12006 0 12042 28 4 br_0_18
port 415 nsew
rlabel metal1 s 12222 0 12258 28 4 br_1_18
port 417 nsew
rlabel metal1 s 12990 0 13026 28 4 bl_0_19
port 419 nsew
rlabel metal1 s 12774 0 12810 28 4 bl_1_19
port 421 nsew
rlabel metal1 s 12918 0 12954 28 4 br_0_19
port 423 nsew
rlabel metal1 s 12702 0 12738 28 4 br_1_19
port 425 nsew
rlabel metal1 s 13182 0 13218 28 4 bl_0_20
port 427 nsew
rlabel metal1 s 13398 0 13434 28 4 bl_1_20
port 429 nsew
rlabel metal1 s 13254 0 13290 28 4 br_0_20
port 431 nsew
rlabel metal1 s 13470 0 13506 28 4 br_1_20
port 433 nsew
rlabel metal1 s 14238 0 14274 28 4 bl_0_21
port 435 nsew
rlabel metal1 s 14022 0 14058 28 4 bl_1_21
port 437 nsew
rlabel metal1 s 14166 0 14202 28 4 br_0_21
port 439 nsew
rlabel metal1 s 13950 0 13986 28 4 br_1_21
port 441 nsew
rlabel metal1 s 14430 0 14466 28 4 bl_0_22
port 443 nsew
rlabel metal1 s 14646 0 14682 28 4 bl_1_22
port 445 nsew
rlabel metal1 s 14502 0 14538 28 4 br_0_22
port 447 nsew
rlabel metal1 s 14718 0 14754 28 4 br_1_22
port 449 nsew
rlabel metal1 s 15486 0 15522 28 4 bl_0_23
port 451 nsew
rlabel metal1 s 15270 0 15306 28 4 bl_1_23
port 453 nsew
rlabel metal1 s 15414 0 15450 28 4 br_0_23
port 455 nsew
rlabel metal1 s 15198 0 15234 28 4 br_1_23
port 457 nsew
rlabel metal1 s 15678 0 15714 28 4 bl_0_24
port 459 nsew
rlabel metal1 s 15894 0 15930 28 4 bl_1_24
port 461 nsew
rlabel metal1 s 15750 0 15786 28 4 br_0_24
port 463 nsew
rlabel metal1 s 15966 0 16002 28 4 br_1_24
port 465 nsew
rlabel metal1 s 16734 0 16770 28 4 bl_0_25
port 467 nsew
rlabel metal1 s 16518 0 16554 28 4 bl_1_25
port 469 nsew
rlabel metal1 s 16662 0 16698 28 4 br_0_25
port 471 nsew
rlabel metal1 s 16446 0 16482 28 4 br_1_25
port 473 nsew
rlabel metal1 s 16926 0 16962 28 4 bl_0_26
port 475 nsew
rlabel metal1 s 17142 0 17178 28 4 bl_1_26
port 477 nsew
rlabel metal1 s 16998 0 17034 28 4 br_0_26
port 479 nsew
rlabel metal1 s 17214 0 17250 28 4 br_1_26
port 481 nsew
rlabel metal1 s 17982 0 18018 28 4 bl_0_27
port 483 nsew
rlabel metal1 s 17766 0 17802 28 4 bl_1_27
port 485 nsew
rlabel metal1 s 17910 0 17946 28 4 br_0_27
port 487 nsew
rlabel metal1 s 17694 0 17730 28 4 br_1_27
port 489 nsew
rlabel metal1 s 18174 0 18210 28 4 bl_0_28
port 491 nsew
rlabel metal1 s 18390 0 18426 28 4 bl_1_28
port 493 nsew
rlabel metal1 s 18246 0 18282 28 4 br_0_28
port 495 nsew
rlabel metal1 s 18462 0 18498 28 4 br_1_28
port 497 nsew
rlabel metal1 s 19230 0 19266 28 4 bl_0_29
port 499 nsew
rlabel metal1 s 19014 0 19050 28 4 bl_1_29
port 501 nsew
rlabel metal1 s 19158 0 19194 28 4 br_0_29
port 503 nsew
rlabel metal1 s 18942 0 18978 28 4 br_1_29
port 505 nsew
rlabel metal1 s 19422 0 19458 28 4 bl_0_30
port 507 nsew
rlabel metal1 s 19638 0 19674 28 4 bl_1_30
port 509 nsew
rlabel metal1 s 19494 0 19530 28 4 br_0_30
port 511 nsew
rlabel metal1 s 19710 0 19746 28 4 br_1_30
port 513 nsew
rlabel metal1 s 20478 0 20514 28 4 bl_0_31
port 515 nsew
rlabel metal1 s 20262 0 20298 28 4 bl_1_31
port 517 nsew
rlabel metal1 s 20406 0 20442 28 4 br_0_31
port 519 nsew
rlabel metal1 s 20190 0 20226 28 4 br_1_31
port 521 nsew
rlabel metal1 s 510 0 546 28 4 rbl_bl_0_0
port 523 nsew
rlabel metal1 s 294 0 330 28 4 rbl_bl_1_0
port 525 nsew
rlabel metal1 s 438 0 474 28 4 rbl_br_0_0
port 527 nsew
rlabel metal1 s 222 0 258 28 4 rbl_br_1_0
port 529 nsew
rlabel metal1 s 20670 0 20706 28 4 rbl_bl_0_1
port 531 nsew
rlabel metal1 s 20886 0 20922 28 4 rbl_bl_1_1
port 533 nsew
rlabel metal1 s 20742 0 20778 28 4 rbl_br_0_1
port 535 nsew
rlabel metal1 s 20958 0 20994 28 4 rbl_br_1_1
port 537 nsew
rlabel metal1 s 7854 765 7890 1106 4 vdd
port 539 nsew
rlabel metal1 s 4590 14694 4626 15035 4 vdd
port 539 nsew
rlabel metal1 s 8334 9164 8370 9505 4 vdd
port 539 nsew
rlabel metal1 s 20814 23384 20850 23725 4 vdd
port 539 nsew
rlabel metal1 s 15342 15775 15378 16116 4 vdd
port 539 nsew
rlabel metal1 s 10350 3925 10386 4266 4 vdd
port 539 nsew
rlabel metal1 s 14094 6295 14130 6636 4 vdd
port 539 nsew
rlabel metal1 s 9582 18145 9618 18486 4 vdd
port 539 nsew
rlabel metal1 s 10350 2844 10386 3185 4 vdd
port 539 nsew
rlabel metal1 s 15822 1264 15858 1605 4 vdd
port 539 nsew
rlabel metal1 s 15342 13904 15378 14245 4 vdd
port 539 nsew
rlabel metal1 s 15342 16274 15378 16615 4 vdd
port 539 nsew
rlabel metal1 s 5358 20224 5394 20565 4 vdd
port 539 nsew
rlabel metal1 s 12078 25754 12114 26095 4 vdd
port 539 nsew
rlabel metal1 s 14574 12324 14610 12665 4 vdd
port 539 nsew
rlabel metal1 s 10830 22095 10866 22436 4 vdd
port 539 nsew
rlabel metal1 s 5358 22594 5394 22935 4 vdd
port 539 nsew
rlabel metal1 s 16590 2345 16626 2686 4 vdd
port 539 nsew
rlabel metal1 s 14094 16274 14130 16615 4 vdd
port 539 nsew
rlabel metal1 s 17070 6794 17106 7135 4 vdd
port 539 nsew
rlabel metal1 s 4590 16565 4626 16906 4 vdd
port 539 nsew
rlabel metal1 s 4590 15484 4626 15825 4 vdd
port 539 nsew
rlabel metal1 s 8334 11035 8370 11376 4 vdd
port 539 nsew
rlabel metal1 s 3342 13405 3378 13746 4 vdd
port 539 nsew
rlabel metal1 s 846 4424 882 4765 4 vdd
port 539 nsew
rlabel metal1 s 4110 9954 4146 10295 4 vdd
port 539 nsew
rlabel metal1 s 17070 474 17106 815 4 vdd
port 539 nsew
rlabel metal1 s 12846 11534 12882 11875 4 vdd
port 539 nsew
rlabel metal1 s 20814 13114 20850 13455 4 vdd
port 539 nsew
rlabel metal1 s 2862 8374 2898 8715 4 vdd
port 539 nsew
rlabel metal1 s 10350 21014 10386 21355 4 vdd
port 539 nsew
rlabel metal1 s 17070 10744 17106 11085 4 vdd
port 539 nsew
rlabel metal1 s 12078 15775 12114 16116 4 vdd
port 539 nsew
rlabel metal1 s 19566 12615 19602 12956 4 vdd
port 539 nsew
rlabel metal1 s 14574 12615 14610 12956 4 vdd
port 539 nsew
rlabel metal1 s 15822 18935 15858 19276 4 vdd
port 539 nsew
rlabel metal1 s 17070 9455 17106 9796 4 vdd
port 539 nsew
rlabel metal1 s 7086 19725 7122 20066 4 vdd
port 539 nsew
rlabel metal1 s 1614 474 1650 815 4 vdd
port 539 nsew
rlabel metal1 s 8334 21804 8370 22145 4 vdd
port 539 nsew
rlabel metal1 s 7086 9164 7122 9505 4 vdd
port 539 nsew
rlabel metal1 s 4110 19434 4146 19775 4 vdd
port 539 nsew
rlabel metal1 s 16590 13904 16626 14245 4 vdd
port 539 nsew
rlabel metal1 s 19086 10744 19122 11085 4 vdd
port 539 nsew
rlabel metal1 s 18318 765 18354 1106 4 vdd
port 539 nsew
rlabel metal1 s 12078 20224 12114 20565 4 vdd
port 539 nsew
rlabel metal1 s 18318 24465 18354 24806 4 vdd
port 539 nsew
rlabel metal1 s 12846 2844 12882 3185 4 vdd
port 539 nsew
rlabel metal1 s 15822 20515 15858 20856 4 vdd
port 539 nsew
rlabel metal1 s 16590 6004 16626 6345 4 vdd
port 539 nsew
rlabel metal1 s 10830 11035 10866 11376 4 vdd
port 539 nsew
rlabel metal1 s 4110 25754 4146 26095 4 vdd
port 539 nsew
rlabel metal1 s 15822 4424 15858 4765 4 vdd
port 539 nsew
rlabel metal1 s 15822 15484 15858 15825 4 vdd
port 539 nsew
rlabel metal1 s 3342 14694 3378 15035 4 vdd
port 539 nsew
rlabel metal1 s 3342 5214 3378 5555 4 vdd
port 539 nsew
rlabel metal1 s 7086 -25 7122 316 4 vdd
port 539 nsew
rlabel metal1 s 11598 14694 11634 15035 4 vdd
port 539 nsew
rlabel metal1 s 2862 7085 2898 7426 4 vdd
port 539 nsew
rlabel metal1 s 11598 6004 11634 6345 4 vdd
port 539 nsew
rlabel metal1 s 20814 9954 20850 10295 4 vdd
port 539 nsew
rlabel metal1 s 14574 9164 14610 9505 4 vdd
port 539 nsew
rlabel metal1 s 20334 24174 20370 24515 4 vdd
port 539 nsew
rlabel metal1 s 9582 9455 9618 9796 4 vdd
port 539 nsew
rlabel metal1 s 11598 11825 11634 12166 4 vdd
port 539 nsew
rlabel metal1 s 17838 -25 17874 316 4 vdd
port 539 nsew
rlabel metal1 s 13326 12615 13362 12956 4 vdd
port 539 nsew
rlabel metal1 s 3342 19725 3378 20066 4 vdd
port 539 nsew
rlabel metal1 s 14094 5505 14130 5846 4 vdd
port 539 nsew
rlabel metal1 s 10830 3135 10866 3476 4 vdd
port 539 nsew
rlabel metal1 s 4110 11825 4146 12166 4 vdd
port 539 nsew
rlabel metal1 s 5358 2345 5394 2686 4 vdd
port 539 nsew
rlabel metal1 s 7086 21014 7122 21355 4 vdd
port 539 nsew
rlabel metal1 s 4590 7584 4626 7925 4 vdd
port 539 nsew
rlabel metal1 s 2862 14195 2898 14536 4 vdd
port 539 nsew
rlabel metal1 s 7086 474 7122 815 4 vdd
port 539 nsew
rlabel metal1 s 5838 3135 5874 3476 4 vdd
port 539 nsew
rlabel metal1 s 17838 13405 17874 13746 4 vdd
port 539 nsew
rlabel metal1 s 15342 18145 15378 18486 4 vdd
port 539 nsew
rlabel metal1 s 19566 14694 19602 15035 4 vdd
port 539 nsew
rlabel metal1 s 13326 25255 13362 25596 4 vdd
port 539 nsew
rlabel metal1 s 4590 2844 4626 3185 4 vdd
port 539 nsew
rlabel metal1 s 15342 9164 15378 9505 4 vdd
port 539 nsew
rlabel metal1 s 5358 7584 5394 7925 4 vdd
port 539 nsew
rlabel metal1 s 15822 19725 15858 20066 4 vdd
port 539 nsew
rlabel metal1 s 3342 8665 3378 9006 4 vdd
port 539 nsew
rlabel metal1 s 3342 8374 3378 8715 4 vdd
port 539 nsew
rlabel metal1 s 10350 1555 10386 1896 4 vdd
port 539 nsew
rlabel metal1 s 2094 19434 2130 19775 4 vdd
port 539 nsew
rlabel metal1 s 9582 24465 9618 24806 4 vdd
port 539 nsew
rlabel metal1 s 5358 20515 5394 20856 4 vdd
port 539 nsew
rlabel metal1 s 17070 17355 17106 17696 4 vdd
port 539 nsew
rlabel metal1 s 1614 8374 1650 8715 4 vdd
port 539 nsew
rlabel metal1 s 14094 18935 14130 19276 4 vdd
port 539 nsew
rlabel metal1 s 20334 6004 20370 6345 4 vdd
port 539 nsew
rlabel metal1 s 846 24465 882 24806 4 vdd
port 539 nsew
rlabel metal1 s 1614 3925 1650 4266 4 vdd
port 539 nsew
rlabel metal1 s 13326 11534 13362 11875 4 vdd
port 539 nsew
rlabel metal1 s 20814 3925 20850 4266 4 vdd
port 539 nsew
rlabel metal1 s 11598 13405 11634 13746 4 vdd
port 539 nsew
rlabel metal1 s 20334 22885 20370 23226 4 vdd
port 539 nsew
rlabel metal1 s 2862 18145 2898 18486 4 vdd
port 539 nsew
rlabel metal1 s 4110 17064 4146 17405 4 vdd
port 539 nsew
rlabel metal1 s 18318 17854 18354 18195 4 vdd
port 539 nsew
rlabel metal1 s 7854 23675 7890 24016 4 vdd
port 539 nsew
rlabel metal1 s 14094 22594 14130 22935 4 vdd
port 539 nsew
rlabel metal1 s 4110 4715 4146 5056 4 vdd
port 539 nsew
rlabel metal1 s 9102 21804 9138 22145 4 vdd
port 539 nsew
rlabel metal1 s 19566 474 19602 815 4 vdd
port 539 nsew
rlabel metal1 s 10350 12615 10386 12956 4 vdd
port 539 nsew
rlabel metal1 s 2094 14985 2130 15326 4 vdd
port 539 nsew
rlabel metal1 s 2862 25754 2898 26095 4 vdd
port 539 nsew
rlabel metal1 s 8334 2054 8370 2395 4 vdd
port 539 nsew
rlabel metal1 s 4110 24964 4146 25305 4 vdd
port 539 nsew
rlabel metal1 s 366 4424 402 4765 4 vdd
port 539 nsew
rlabel metal1 s 6606 474 6642 815 4 vdd
port 539 nsew
rlabel metal1 s 9582 1264 9618 1605 4 vdd
port 539 nsew
rlabel metal1 s 3342 3925 3378 4266 4 vdd
port 539 nsew
rlabel metal1 s 4590 -25 4626 316 4 vdd
port 539 nsew
rlabel metal1 s 6606 7085 6642 7426 4 vdd
port 539 nsew
rlabel metal1 s 17070 17854 17106 18195 4 vdd
port 539 nsew
rlabel metal1 s 18318 17064 18354 17405 4 vdd
port 539 nsew
rlabel metal1 s 6606 5214 6642 5555 4 vdd
port 539 nsew
rlabel metal1 s 13326 6004 13362 6345 4 vdd
port 539 nsew
rlabel metal1 s 12078 13405 12114 13746 4 vdd
port 539 nsew
rlabel metal1 s 13326 24465 13362 24806 4 vdd
port 539 nsew
rlabel metal1 s 20814 2054 20850 2395 4 vdd
port 539 nsew
rlabel metal1 s 7086 7584 7122 7925 4 vdd
port 539 nsew
rlabel metal1 s 10830 2345 10866 2686 4 vdd
port 539 nsew
rlabel metal1 s 19086 13114 19122 13455 4 vdd
port 539 nsew
rlabel metal1 s 9582 8665 9618 9006 4 vdd
port 539 nsew
rlabel metal1 s 2862 11035 2898 11376 4 vdd
port 539 nsew
rlabel metal1 s 10830 21014 10866 21355 4 vdd
port 539 nsew
rlabel metal1 s 9102 16274 9138 16615 4 vdd
port 539 nsew
rlabel metal1 s 4110 -25 4146 316 4 vdd
port 539 nsew
rlabel metal1 s 4590 9954 4626 10295 4 vdd
port 539 nsew
rlabel metal1 s 8334 5214 8370 5555 4 vdd
port 539 nsew
rlabel metal1 s 7086 6295 7122 6636 4 vdd
port 539 nsew
rlabel metal1 s 4110 12615 4146 12956 4 vdd
port 539 nsew
rlabel metal1 s 17070 14985 17106 15326 4 vdd
port 539 nsew
rlabel metal1 s 11598 3135 11634 3476 4 vdd
port 539 nsew
rlabel metal1 s 5358 14195 5394 14536 4 vdd
port 539 nsew
rlabel metal1 s 9582 15484 9618 15825 4 vdd
port 539 nsew
rlabel metal1 s 15822 4715 15858 5056 4 vdd
port 539 nsew
rlabel metal1 s 846 22095 882 22436 4 vdd
port 539 nsew
rlabel metal1 s 14094 7085 14130 7426 4 vdd
port 539 nsew
rlabel metal1 s 20334 16565 20370 16906 4 vdd
port 539 nsew
rlabel metal1 s 5358 23675 5394 24016 4 vdd
port 539 nsew
rlabel metal1 s 4110 13114 4146 13455 4 vdd
port 539 nsew
rlabel metal1 s 17070 19434 17106 19775 4 vdd
port 539 nsew
rlabel metal1 s 7086 2054 7122 2395 4 vdd
port 539 nsew
rlabel metal1 s 366 7085 402 7426 4 vdd
port 539 nsew
rlabel metal1 s 366 19725 402 20066 4 vdd
port 539 nsew
rlabel metal1 s 9582 16274 9618 16615 4 vdd
port 539 nsew
rlabel metal1 s 12078 2054 12114 2395 4 vdd
port 539 nsew
rlabel metal1 s 17838 9164 17874 9505 4 vdd
port 539 nsew
rlabel metal1 s 16590 13405 16626 13746 4 vdd
port 539 nsew
rlabel metal1 s 8334 7085 8370 7426 4 vdd
port 539 nsew
rlabel metal1 s 16590 20224 16626 20565 4 vdd
port 539 nsew
rlabel metal1 s 5358 9164 5394 9505 4 vdd
port 539 nsew
rlabel metal1 s 2094 22885 2130 23226 4 vdd
port 539 nsew
rlabel metal1 s 4110 10744 4146 11085 4 vdd
port 539 nsew
rlabel metal1 s 18318 23675 18354 24016 4 vdd
port 539 nsew
rlabel metal1 s 4590 4715 4626 5056 4 vdd
port 539 nsew
rlabel metal1 s 1614 24174 1650 24515 4 vdd
port 539 nsew
rlabel metal1 s 18318 3634 18354 3975 4 vdd
port 539 nsew
rlabel metal1 s 11598 13904 11634 14245 4 vdd
port 539 nsew
rlabel metal1 s 13326 4715 13362 5056 4 vdd
port 539 nsew
rlabel metal1 s 12078 3634 12114 3975 4 vdd
port 539 nsew
rlabel metal1 s 10350 19434 10386 19775 4 vdd
port 539 nsew
rlabel metal1 s 13326 765 13362 1106 4 vdd
port 539 nsew
rlabel metal1 s 11598 22095 11634 22436 4 vdd
port 539 nsew
rlabel metal1 s 366 20224 402 20565 4 vdd
port 539 nsew
rlabel metal1 s 20814 21804 20850 22145 4 vdd
port 539 nsew
rlabel metal1 s 17070 14694 17106 15035 4 vdd
port 539 nsew
rlabel metal1 s 2094 2345 2130 2686 4 vdd
port 539 nsew
rlabel metal1 s 17838 20515 17874 20856 4 vdd
port 539 nsew
rlabel metal1 s 7854 10245 7890 10586 4 vdd
port 539 nsew
rlabel metal1 s 12078 7085 12114 7426 4 vdd
port 539 nsew
rlabel metal1 s 17070 6295 17106 6636 4 vdd
port 539 nsew
rlabel metal1 s 9582 21305 9618 21646 4 vdd
port 539 nsew
rlabel metal1 s 4110 14694 4146 15035 4 vdd
port 539 nsew
rlabel metal1 s 15822 3925 15858 4266 4 vdd
port 539 nsew
rlabel metal1 s 6606 2054 6642 2395 4 vdd
port 539 nsew
rlabel metal1 s 6606 3925 6642 4266 4 vdd
port 539 nsew
rlabel metal1 s 12846 20224 12882 20565 4 vdd
port 539 nsew
rlabel metal1 s 20814 23675 20850 24016 4 vdd
port 539 nsew
rlabel metal1 s 19566 16274 19602 16615 4 vdd
port 539 nsew
rlabel metal1 s 7854 22885 7890 23226 4 vdd
port 539 nsew
rlabel metal1 s 9582 19434 9618 19775 4 vdd
port 539 nsew
rlabel metal1 s 7086 9455 7122 9796 4 vdd
port 539 nsew
rlabel metal1 s 4110 1555 4146 1896 4 vdd
port 539 nsew
rlabel metal1 s 14094 23675 14130 24016 4 vdd
port 539 nsew
rlabel metal1 s 19086 15775 19122 16116 4 vdd
port 539 nsew
rlabel metal1 s 15822 24174 15858 24515 4 vdd
port 539 nsew
rlabel metal1 s 12078 2345 12114 2686 4 vdd
port 539 nsew
rlabel metal1 s 13326 2345 13362 2686 4 vdd
port 539 nsew
rlabel metal1 s 14574 11035 14610 11376 4 vdd
port 539 nsew
rlabel metal1 s 5358 11825 5394 12166 4 vdd
port 539 nsew
rlabel metal1 s 2094 6004 2130 6345 4 vdd
port 539 nsew
rlabel metal1 s 10830 23675 10866 24016 4 vdd
port 539 nsew
rlabel metal1 s 19566 18644 19602 18985 4 vdd
port 539 nsew
rlabel metal1 s 14094 11035 14130 11376 4 vdd
port 539 nsew
rlabel metal1 s 12846 16565 12882 16906 4 vdd
port 539 nsew
rlabel metal1 s 15822 765 15858 1106 4 vdd
port 539 nsew
rlabel metal1 s 18318 4715 18354 5056 4 vdd
port 539 nsew
rlabel metal1 s 15342 17355 15378 17696 4 vdd
port 539 nsew
rlabel metal1 s 19086 18644 19122 18985 4 vdd
port 539 nsew
rlabel metal1 s 2862 6794 2898 7135 4 vdd
port 539 nsew
rlabel metal1 s 20334 9954 20370 10295 4 vdd
port 539 nsew
rlabel metal1 s 5838 3634 5874 3975 4 vdd
port 539 nsew
rlabel metal1 s 2862 1264 2898 1605 4 vdd
port 539 nsew
rlabel metal1 s 5358 5505 5394 5846 4 vdd
port 539 nsew
rlabel metal1 s 12078 6794 12114 7135 4 vdd
port 539 nsew
rlabel metal1 s 2862 17854 2898 18195 4 vdd
port 539 nsew
rlabel metal1 s 14574 14985 14610 15326 4 vdd
port 539 nsew
rlabel metal1 s 17070 21305 17106 21646 4 vdd
port 539 nsew
rlabel metal1 s 15342 19725 15378 20066 4 vdd
port 539 nsew
rlabel metal1 s 12846 9954 12882 10295 4 vdd
port 539 nsew
rlabel metal1 s 12846 18935 12882 19276 4 vdd
port 539 nsew
rlabel metal1 s 16590 2054 16626 2395 4 vdd
port 539 nsew
rlabel metal1 s 13326 23384 13362 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 16565 8370 16906 4 vdd
port 539 nsew
rlabel metal1 s 17838 4715 17874 5056 4 vdd
port 539 nsew
rlabel metal1 s 16590 7085 16626 7426 4 vdd
port 539 nsew
rlabel metal1 s 13326 8665 13362 9006 4 vdd
port 539 nsew
rlabel metal1 s 18318 15484 18354 15825 4 vdd
port 539 nsew
rlabel metal1 s 16590 11035 16626 11376 4 vdd
port 539 nsew
rlabel metal1 s 846 17064 882 17405 4 vdd
port 539 nsew
rlabel metal1 s 16590 25754 16626 26095 4 vdd
port 539 nsew
rlabel metal1 s 20814 6794 20850 7135 4 vdd
port 539 nsew
rlabel metal1 s 12846 3634 12882 3975 4 vdd
port 539 nsew
rlabel metal1 s 12846 21305 12882 21646 4 vdd
port 539 nsew
rlabel metal1 s 12846 14694 12882 15035 4 vdd
port 539 nsew
rlabel metal1 s 4590 8374 4626 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 7085 9138 7426 4 vdd
port 539 nsew
rlabel metal1 s 17070 7085 17106 7426 4 vdd
port 539 nsew
rlabel metal1 s 19566 6295 19602 6636 4 vdd
port 539 nsew
rlabel metal1 s 1614 18145 1650 18486 4 vdd
port 539 nsew
rlabel metal1 s 14094 25754 14130 26095 4 vdd
port 539 nsew
rlabel metal1 s 12846 23675 12882 24016 4 vdd
port 539 nsew
rlabel metal1 s 18318 14195 18354 14536 4 vdd
port 539 nsew
rlabel metal1 s 5838 7875 5874 8216 4 vdd
port 539 nsew
rlabel metal1 s 14574 25255 14610 25596 4 vdd
port 539 nsew
rlabel metal1 s 7086 17064 7122 17405 4 vdd
port 539 nsew
rlabel metal1 s 1614 6794 1650 7135 4 vdd
port 539 nsew
rlabel metal1 s 3342 7085 3378 7426 4 vdd
port 539 nsew
rlabel metal1 s 12078 14985 12114 15326 4 vdd
port 539 nsew
rlabel metal1 s 10350 24174 10386 24515 4 vdd
port 539 nsew
rlabel metal1 s 9582 12615 9618 12956 4 vdd
port 539 nsew
rlabel metal1 s 846 17355 882 17696 4 vdd
port 539 nsew
rlabel metal1 s 9582 2054 9618 2395 4 vdd
port 539 nsew
rlabel metal1 s 4590 20515 4626 20856 4 vdd
port 539 nsew
rlabel metal1 s 4590 14985 4626 15326 4 vdd
port 539 nsew
rlabel metal1 s 7854 9954 7890 10295 4 vdd
port 539 nsew
rlabel metal1 s 846 11825 882 12166 4 vdd
port 539 nsew
rlabel metal1 s 2094 23384 2130 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 21305 8370 21646 4 vdd
port 539 nsew
rlabel metal1 s 366 21305 402 21646 4 vdd
port 539 nsew
rlabel metal1 s 17070 18935 17106 19276 4 vdd
port 539 nsew
rlabel metal1 s 15822 17064 15858 17405 4 vdd
port 539 nsew
rlabel metal1 s 2094 17064 2130 17405 4 vdd
port 539 nsew
rlabel metal1 s 9102 2844 9138 3185 4 vdd
port 539 nsew
rlabel metal1 s 5838 22095 5874 22436 4 vdd
port 539 nsew
rlabel metal1 s 18318 3925 18354 4266 4 vdd
port 539 nsew
rlabel metal1 s 7086 21804 7122 22145 4 vdd
port 539 nsew
rlabel metal1 s 9582 17064 9618 17405 4 vdd
port 539 nsew
rlabel metal1 s 1614 22594 1650 22935 4 vdd
port 539 nsew
rlabel metal1 s 7086 22885 7122 23226 4 vdd
port 539 nsew
rlabel metal1 s 1614 3135 1650 3476 4 vdd
port 539 nsew
rlabel metal1 s 8334 2844 8370 3185 4 vdd
port 539 nsew
rlabel metal1 s 9102 21014 9138 21355 4 vdd
port 539 nsew
rlabel metal1 s 12846 22095 12882 22436 4 vdd
port 539 nsew
rlabel metal1 s 7086 16565 7122 16906 4 vdd
port 539 nsew
rlabel metal1 s 15342 12615 15378 12956 4 vdd
port 539 nsew
rlabel metal1 s 12846 22885 12882 23226 4 vdd
port 539 nsew
rlabel metal1 s 5838 16274 5874 16615 4 vdd
port 539 nsew
rlabel metal1 s 5358 25255 5394 25596 4 vdd
port 539 nsew
rlabel metal1 s 14574 -25 14610 316 4 vdd
port 539 nsew
rlabel metal1 s 18318 18644 18354 18985 4 vdd
port 539 nsew
rlabel metal1 s 1614 9164 1650 9505 4 vdd
port 539 nsew
rlabel metal1 s 17838 18935 17874 19276 4 vdd
port 539 nsew
rlabel metal1 s 13326 18145 13362 18486 4 vdd
port 539 nsew
rlabel metal1 s 8334 11825 8370 12166 4 vdd
port 539 nsew
rlabel metal1 s 17070 20515 17106 20856 4 vdd
port 539 nsew
rlabel metal1 s 17838 16565 17874 16906 4 vdd
port 539 nsew
rlabel metal1 s 4110 13405 4146 13746 4 vdd
port 539 nsew
rlabel metal1 s 10830 23384 10866 23725 4 vdd
port 539 nsew
rlabel metal1 s 10830 25255 10866 25596 4 vdd
port 539 nsew
rlabel metal1 s 12846 7085 12882 7426 4 vdd
port 539 nsew
rlabel metal1 s 10350 13904 10386 14245 4 vdd
port 539 nsew
rlabel metal1 s 9102 5505 9138 5846 4 vdd
port 539 nsew
rlabel metal1 s 12078 5505 12114 5846 4 vdd
port 539 nsew
rlabel metal1 s 4110 18644 4146 18985 4 vdd
port 539 nsew
rlabel metal1 s 10830 6004 10866 6345 4 vdd
port 539 nsew
rlabel metal1 s 10830 12615 10866 12956 4 vdd
port 539 nsew
rlabel metal1 s 3342 2345 3378 2686 4 vdd
port 539 nsew
rlabel metal1 s 10830 765 10866 1106 4 vdd
port 539 nsew
rlabel metal1 s 2094 10744 2130 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 3925 14610 4266 4 vdd
port 539 nsew
rlabel metal1 s 16590 3925 16626 4266 4 vdd
port 539 nsew
rlabel metal1 s 366 17355 402 17696 4 vdd
port 539 nsew
rlabel metal1 s 15342 10245 15378 10586 4 vdd
port 539 nsew
rlabel metal1 s 17838 17854 17874 18195 4 vdd
port 539 nsew
rlabel metal1 s 14574 17064 14610 17405 4 vdd
port 539 nsew
rlabel metal1 s 17838 5214 17874 5555 4 vdd
port 539 nsew
rlabel metal1 s 11598 18935 11634 19276 4 vdd
port 539 nsew
rlabel metal1 s 20814 9455 20850 9796 4 vdd
port 539 nsew
rlabel metal1 s 846 14195 882 14536 4 vdd
port 539 nsew
rlabel metal1 s 1614 21014 1650 21355 4 vdd
port 539 nsew
rlabel metal1 s 12078 17854 12114 18195 4 vdd
port 539 nsew
rlabel metal1 s 7854 2054 7890 2395 4 vdd
port 539 nsew
rlabel metal1 s 9582 17355 9618 17696 4 vdd
port 539 nsew
rlabel metal1 s 2862 18935 2898 19276 4 vdd
port 539 nsew
rlabel metal1 s 17838 11035 17874 11376 4 vdd
port 539 nsew
rlabel metal1 s 9582 6794 9618 7135 4 vdd
port 539 nsew
rlabel metal1 s 4110 9455 4146 9796 4 vdd
port 539 nsew
rlabel metal1 s 5838 21804 5874 22145 4 vdd
port 539 nsew
rlabel metal1 s 9582 14195 9618 14536 4 vdd
port 539 nsew
rlabel metal1 s 6606 25255 6642 25596 4 vdd
port 539 nsew
rlabel metal1 s 20334 20515 20370 20856 4 vdd
port 539 nsew
rlabel metal1 s 6606 24964 6642 25305 4 vdd
port 539 nsew
rlabel metal1 s 15342 8665 15378 9006 4 vdd
port 539 nsew
rlabel metal1 s 2094 19725 2130 20066 4 vdd
port 539 nsew
rlabel metal1 s 18318 19725 18354 20066 4 vdd
port 539 nsew
rlabel metal1 s 846 12324 882 12665 4 vdd
port 539 nsew
rlabel metal1 s 2862 14694 2898 15035 4 vdd
port 539 nsew
rlabel metal1 s 18318 23384 18354 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 11534 8370 11875 4 vdd
port 539 nsew
rlabel metal1 s 17070 22594 17106 22935 4 vdd
port 539 nsew
rlabel metal1 s 17070 10245 17106 10586 4 vdd
port 539 nsew
rlabel metal1 s 7854 11035 7890 11376 4 vdd
port 539 nsew
rlabel metal1 s 2862 15484 2898 15825 4 vdd
port 539 nsew
rlabel metal1 s 14574 11825 14610 12166 4 vdd
port 539 nsew
rlabel metal1 s 5358 13405 5394 13746 4 vdd
port 539 nsew
rlabel metal1 s 18318 7085 18354 7426 4 vdd
port 539 nsew
rlabel metal1 s 13326 3925 13362 4266 4 vdd
port 539 nsew
rlabel metal1 s 19566 25255 19602 25596 4 vdd
port 539 nsew
rlabel metal1 s 10830 15775 10866 16116 4 vdd
port 539 nsew
rlabel metal1 s 7854 5214 7890 5555 4 vdd
port 539 nsew
rlabel metal1 s 11598 12324 11634 12665 4 vdd
port 539 nsew
rlabel metal1 s 5358 1555 5394 1896 4 vdd
port 539 nsew
rlabel metal1 s 11598 25754 11634 26095 4 vdd
port 539 nsew
rlabel metal1 s 3342 10245 3378 10586 4 vdd
port 539 nsew
rlabel metal1 s 11598 16565 11634 16906 4 vdd
port 539 nsew
rlabel metal1 s 13326 25754 13362 26095 4 vdd
port 539 nsew
rlabel metal1 s 14094 4715 14130 5056 4 vdd
port 539 nsew
rlabel metal1 s 846 24174 882 24515 4 vdd
port 539 nsew
rlabel metal1 s 1614 7085 1650 7426 4 vdd
port 539 nsew
rlabel metal1 s 15342 21804 15378 22145 4 vdd
port 539 nsew
rlabel metal1 s 18318 5214 18354 5555 4 vdd
port 539 nsew
rlabel metal1 s 14094 13904 14130 14245 4 vdd
port 539 nsew
rlabel metal1 s 846 13405 882 13746 4 vdd
port 539 nsew
rlabel metal1 s 19566 21305 19602 21646 4 vdd
port 539 nsew
rlabel metal1 s 19086 24964 19122 25305 4 vdd
port 539 nsew
rlabel metal1 s 12846 6295 12882 6636 4 vdd
port 539 nsew
rlabel metal1 s 11598 21305 11634 21646 4 vdd
port 539 nsew
rlabel metal1 s 846 16565 882 16906 4 vdd
port 539 nsew
rlabel metal1 s 1614 10744 1650 11085 4 vdd
port 539 nsew
rlabel metal1 s 366 3634 402 3975 4 vdd
port 539 nsew
rlabel metal1 s 15342 4715 15378 5056 4 vdd
port 539 nsew
rlabel metal1 s 14574 5214 14610 5555 4 vdd
port 539 nsew
rlabel metal1 s 5838 7085 5874 7426 4 vdd
port 539 nsew
rlabel metal1 s 12078 21014 12114 21355 4 vdd
port 539 nsew
rlabel metal1 s 366 22885 402 23226 4 vdd
port 539 nsew
rlabel metal1 s 17070 11035 17106 11376 4 vdd
port 539 nsew
rlabel metal1 s 12846 765 12882 1106 4 vdd
port 539 nsew
rlabel metal1 s 14094 15484 14130 15825 4 vdd
port 539 nsew
rlabel metal1 s 15822 -25 15858 316 4 vdd
port 539 nsew
rlabel metal1 s 9582 3135 9618 3476 4 vdd
port 539 nsew
rlabel metal1 s 366 474 402 815 4 vdd
port 539 nsew
rlabel metal1 s 20814 10744 20850 11085 4 vdd
port 539 nsew
rlabel metal1 s 4590 23675 4626 24016 4 vdd
port 539 nsew
rlabel metal1 s 2862 10245 2898 10586 4 vdd
port 539 nsew
rlabel metal1 s 2094 24174 2130 24515 4 vdd
port 539 nsew
rlabel metal1 s 5358 18145 5394 18486 4 vdd
port 539 nsew
rlabel metal1 s 8334 15484 8370 15825 4 vdd
port 539 nsew
rlabel metal1 s 5358 24465 5394 24806 4 vdd
port 539 nsew
rlabel metal1 s 14094 22885 14130 23226 4 vdd
port 539 nsew
rlabel metal1 s 5838 6295 5874 6636 4 vdd
port 539 nsew
rlabel metal1 s 17838 3634 17874 3975 4 vdd
port 539 nsew
rlabel metal1 s 4110 22095 4146 22436 4 vdd
port 539 nsew
rlabel metal1 s 366 13904 402 14245 4 vdd
port 539 nsew
rlabel metal1 s 15342 9954 15378 10295 4 vdd
port 539 nsew
rlabel metal1 s 9102 14195 9138 14536 4 vdd
port 539 nsew
rlabel metal1 s 7086 8374 7122 8715 4 vdd
port 539 nsew
rlabel metal1 s 5838 18935 5874 19276 4 vdd
port 539 nsew
rlabel metal1 s 16590 1555 16626 1896 4 vdd
port 539 nsew
rlabel metal1 s 7854 24174 7890 24515 4 vdd
port 539 nsew
rlabel metal1 s 11598 5214 11634 5555 4 vdd
port 539 nsew
rlabel metal1 s 16590 19434 16626 19775 4 vdd
port 539 nsew
rlabel metal1 s 12078 22594 12114 22935 4 vdd
port 539 nsew
rlabel metal1 s 7854 16565 7890 16906 4 vdd
port 539 nsew
rlabel metal1 s 12846 11825 12882 12166 4 vdd
port 539 nsew
rlabel metal1 s 4590 23384 4626 23725 4 vdd
port 539 nsew
rlabel metal1 s 2094 7875 2130 8216 4 vdd
port 539 nsew
rlabel metal1 s 10350 2054 10386 2395 4 vdd
port 539 nsew
rlabel metal1 s 6606 21804 6642 22145 4 vdd
port 539 nsew
rlabel metal1 s 6606 18644 6642 18985 4 vdd
port 539 nsew
rlabel metal1 s 15342 24964 15378 25305 4 vdd
port 539 nsew
rlabel metal1 s 8334 25754 8370 26095 4 vdd
port 539 nsew
rlabel metal1 s 10830 1264 10866 1605 4 vdd
port 539 nsew
rlabel metal1 s 8334 10744 8370 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 2345 14610 2686 4 vdd
port 539 nsew
rlabel metal1 s 11598 17854 11634 18195 4 vdd
port 539 nsew
rlabel metal1 s 5358 11035 5394 11376 4 vdd
port 539 nsew
rlabel metal1 s 20814 22095 20850 22436 4 vdd
port 539 nsew
rlabel metal1 s 15342 474 15378 815 4 vdd
port 539 nsew
rlabel metal1 s 5358 13904 5394 14245 4 vdd
port 539 nsew
rlabel metal1 s 10350 7584 10386 7925 4 vdd
port 539 nsew
rlabel metal1 s 7086 16274 7122 16615 4 vdd
port 539 nsew
rlabel metal1 s 4590 21305 4626 21646 4 vdd
port 539 nsew
rlabel metal1 s 2094 13904 2130 14245 4 vdd
port 539 nsew
rlabel metal1 s 11598 13114 11634 13455 4 vdd
port 539 nsew
rlabel metal1 s 16590 11825 16626 12166 4 vdd
port 539 nsew
rlabel metal1 s 20814 17854 20850 18195 4 vdd
port 539 nsew
rlabel metal1 s 12078 21305 12114 21646 4 vdd
port 539 nsew
rlabel metal1 s 8334 17355 8370 17696 4 vdd
port 539 nsew
rlabel metal1 s 846 4715 882 5056 4 vdd
port 539 nsew
rlabel metal1 s 19566 13114 19602 13455 4 vdd
port 539 nsew
rlabel metal1 s 19566 21014 19602 21355 4 vdd
port 539 nsew
rlabel metal1 s 10350 14985 10386 15326 4 vdd
port 539 nsew
rlabel metal1 s 12846 -25 12882 316 4 vdd
port 539 nsew
rlabel metal1 s 6606 9954 6642 10295 4 vdd
port 539 nsew
rlabel metal1 s 2862 9164 2898 9505 4 vdd
port 539 nsew
rlabel metal1 s 17838 22594 17874 22935 4 vdd
port 539 nsew
rlabel metal1 s 20814 17064 20850 17405 4 vdd
port 539 nsew
rlabel metal1 s 846 7085 882 7426 4 vdd
port 539 nsew
rlabel metal1 s 14574 1555 14610 1896 4 vdd
port 539 nsew
rlabel metal1 s 16590 10245 16626 10586 4 vdd
port 539 nsew
rlabel metal1 s 14094 25255 14130 25596 4 vdd
port 539 nsew
rlabel metal1 s 7086 13904 7122 14245 4 vdd
port 539 nsew
rlabel metal1 s 9582 -25 9618 316 4 vdd
port 539 nsew
rlabel metal1 s 5358 21804 5394 22145 4 vdd
port 539 nsew
rlabel metal1 s 10830 12324 10866 12665 4 vdd
port 539 nsew
rlabel metal1 s 7086 24174 7122 24515 4 vdd
port 539 nsew
rlabel metal1 s 17838 13904 17874 14245 4 vdd
port 539 nsew
rlabel metal1 s 5838 6794 5874 7135 4 vdd
port 539 nsew
rlabel metal1 s 10350 21305 10386 21646 4 vdd
port 539 nsew
rlabel metal1 s 9582 19725 9618 20066 4 vdd
port 539 nsew
rlabel metal1 s 6606 4424 6642 4765 4 vdd
port 539 nsew
rlabel metal1 s 7086 14195 7122 14536 4 vdd
port 539 nsew
rlabel metal1 s 6606 14195 6642 14536 4 vdd
port 539 nsew
rlabel metal1 s 5358 24174 5394 24515 4 vdd
port 539 nsew
rlabel metal1 s 12846 474 12882 815 4 vdd
port 539 nsew
rlabel metal1 s 2862 6295 2898 6636 4 vdd
port 539 nsew
rlabel metal1 s 13326 22885 13362 23226 4 vdd
port 539 nsew
rlabel metal1 s 5838 17854 5874 18195 4 vdd
port 539 nsew
rlabel metal1 s 3342 7584 3378 7925 4 vdd
port 539 nsew
rlabel metal1 s 17838 17355 17874 17696 4 vdd
port 539 nsew
rlabel metal1 s 8334 6295 8370 6636 4 vdd
port 539 nsew
rlabel metal1 s 6606 18935 6642 19276 4 vdd
port 539 nsew
rlabel metal1 s 2862 24174 2898 24515 4 vdd
port 539 nsew
rlabel metal1 s 17070 5505 17106 5846 4 vdd
port 539 nsew
rlabel metal1 s 12846 2345 12882 2686 4 vdd
port 539 nsew
rlabel metal1 s 14574 24964 14610 25305 4 vdd
port 539 nsew
rlabel metal1 s 1614 23384 1650 23725 4 vdd
port 539 nsew
rlabel metal1 s 7854 3135 7890 3476 4 vdd
port 539 nsew
rlabel metal1 s 15822 18644 15858 18985 4 vdd
port 539 nsew
rlabel metal1 s 16590 4424 16626 4765 4 vdd
port 539 nsew
rlabel metal1 s 9102 9954 9138 10295 4 vdd
port 539 nsew
rlabel metal1 s 3342 16565 3378 16906 4 vdd
port 539 nsew
rlabel metal1 s 20814 13405 20850 13746 4 vdd
port 539 nsew
rlabel metal1 s 12078 1555 12114 1896 4 vdd
port 539 nsew
rlabel metal1 s 1614 13114 1650 13455 4 vdd
port 539 nsew
rlabel metal1 s 17838 15484 17874 15825 4 vdd
port 539 nsew
rlabel metal1 s 19566 14985 19602 15326 4 vdd
port 539 nsew
rlabel metal1 s 15342 7085 15378 7426 4 vdd
port 539 nsew
rlabel metal1 s 14094 6004 14130 6345 4 vdd
port 539 nsew
rlabel metal1 s 2862 16274 2898 16615 4 vdd
port 539 nsew
rlabel metal1 s 7086 25255 7122 25596 4 vdd
port 539 nsew
rlabel metal1 s 5838 12324 5874 12665 4 vdd
port 539 nsew
rlabel metal1 s 366 25754 402 26095 4 vdd
port 539 nsew
rlabel metal1 s 10830 8665 10866 9006 4 vdd
port 539 nsew
rlabel metal1 s 6606 8374 6642 8715 4 vdd
port 539 nsew
rlabel metal1 s 20334 8665 20370 9006 4 vdd
port 539 nsew
rlabel metal1 s 16590 3135 16626 3476 4 vdd
port 539 nsew
rlabel metal1 s 20814 11035 20850 11376 4 vdd
port 539 nsew
rlabel metal1 s 14574 765 14610 1106 4 vdd
port 539 nsew
rlabel metal1 s 4110 8665 4146 9006 4 vdd
port 539 nsew
rlabel metal1 s 5358 2844 5394 3185 4 vdd
port 539 nsew
rlabel metal1 s 11598 14195 11634 14536 4 vdd
port 539 nsew
rlabel metal1 s 15342 18644 15378 18985 4 vdd
port 539 nsew
rlabel metal1 s 3342 3634 3378 3975 4 vdd
port 539 nsew
rlabel metal1 s 18318 21014 18354 21355 4 vdd
port 539 nsew
rlabel metal1 s 846 23384 882 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 14694 8370 15035 4 vdd
port 539 nsew
rlabel metal1 s 7086 25754 7122 26095 4 vdd
port 539 nsew
rlabel metal1 s 6606 19725 6642 20066 4 vdd
port 539 nsew
rlabel metal1 s 9582 15775 9618 16116 4 vdd
port 539 nsew
rlabel metal1 s 2862 17355 2898 17696 4 vdd
port 539 nsew
rlabel metal1 s 18318 10744 18354 11085 4 vdd
port 539 nsew
rlabel metal1 s 846 21014 882 21355 4 vdd
port 539 nsew
rlabel metal1 s 9582 22594 9618 22935 4 vdd
port 539 nsew
rlabel metal1 s 366 14985 402 15326 4 vdd
port 539 nsew
rlabel metal1 s 15342 23384 15378 23725 4 vdd
port 539 nsew
rlabel metal1 s 19086 3634 19122 3975 4 vdd
port 539 nsew
rlabel metal1 s 1614 6004 1650 6345 4 vdd
port 539 nsew
rlabel metal1 s 8334 12615 8370 12956 4 vdd
port 539 nsew
rlabel metal1 s 5358 18935 5394 19276 4 vdd
port 539 nsew
rlabel metal1 s 4590 3925 4626 4266 4 vdd
port 539 nsew
rlabel metal1 s 20814 24174 20850 24515 4 vdd
port 539 nsew
rlabel metal1 s 20814 4715 20850 5056 4 vdd
port 539 nsew
rlabel metal1 s 846 21804 882 22145 4 vdd
port 539 nsew
rlabel metal1 s 4590 7085 4626 7426 4 vdd
port 539 nsew
rlabel metal1 s 14094 19434 14130 19775 4 vdd
port 539 nsew
rlabel metal1 s 13326 16274 13362 16615 4 vdd
port 539 nsew
rlabel metal1 s 15342 3135 15378 3476 4 vdd
port 539 nsew
rlabel metal1 s 11598 22594 11634 22935 4 vdd
port 539 nsew
rlabel metal1 s 3342 6295 3378 6636 4 vdd
port 539 nsew
rlabel metal1 s 1614 20224 1650 20565 4 vdd
port 539 nsew
rlabel metal1 s 20814 19434 20850 19775 4 vdd
port 539 nsew
rlabel metal1 s 15822 21014 15858 21355 4 vdd
port 539 nsew
rlabel metal1 s 366 13114 402 13455 4 vdd
port 539 nsew
rlabel metal1 s 18318 8374 18354 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 18145 9138 18486 4 vdd
port 539 nsew
rlabel metal1 s 20334 3135 20370 3476 4 vdd
port 539 nsew
rlabel metal1 s 11598 3634 11634 3975 4 vdd
port 539 nsew
rlabel metal1 s 17070 8665 17106 9006 4 vdd
port 539 nsew
rlabel metal1 s 366 6295 402 6636 4 vdd
port 539 nsew
rlabel metal1 s 13326 1555 13362 1896 4 vdd
port 539 nsew
rlabel metal1 s 3342 21804 3378 22145 4 vdd
port 539 nsew
rlabel metal1 s 4110 16565 4146 16906 4 vdd
port 539 nsew
rlabel metal1 s 20334 21305 20370 21646 4 vdd
port 539 nsew
rlabel metal1 s 17838 12615 17874 12956 4 vdd
port 539 nsew
rlabel metal1 s 3342 4424 3378 4765 4 vdd
port 539 nsew
rlabel metal1 s 17838 14985 17874 15326 4 vdd
port 539 nsew
rlabel metal1 s 17070 24964 17106 25305 4 vdd
port 539 nsew
rlabel metal1 s 14574 1264 14610 1605 4 vdd
port 539 nsew
rlabel metal1 s 17838 14694 17874 15035 4 vdd
port 539 nsew
rlabel metal1 s 6606 14694 6642 15035 4 vdd
port 539 nsew
rlabel metal1 s 5358 17355 5394 17696 4 vdd
port 539 nsew
rlabel metal1 s 12078 16565 12114 16906 4 vdd
port 539 nsew
rlabel metal1 s 12078 9455 12114 9796 4 vdd
port 539 nsew
rlabel metal1 s 2862 765 2898 1106 4 vdd
port 539 nsew
rlabel metal1 s 12846 6794 12882 7135 4 vdd
port 539 nsew
rlabel metal1 s 2094 1555 2130 1896 4 vdd
port 539 nsew
rlabel metal1 s 9582 7584 9618 7925 4 vdd
port 539 nsew
rlabel metal1 s 2862 3135 2898 3476 4 vdd
port 539 nsew
rlabel metal1 s 1614 19434 1650 19775 4 vdd
port 539 nsew
rlabel metal1 s 366 16274 402 16615 4 vdd
port 539 nsew
rlabel metal1 s 1614 13904 1650 14245 4 vdd
port 539 nsew
rlabel metal1 s 2862 22885 2898 23226 4 vdd
port 539 nsew
rlabel metal1 s 12078 -25 12114 316 4 vdd
port 539 nsew
rlabel metal1 s 14574 9455 14610 9796 4 vdd
port 539 nsew
rlabel metal1 s 14574 21804 14610 22145 4 vdd
port 539 nsew
rlabel metal1 s 3342 19434 3378 19775 4 vdd
port 539 nsew
rlabel metal1 s 15822 8665 15858 9006 4 vdd
port 539 nsew
rlabel metal1 s 10830 13114 10866 13455 4 vdd
port 539 nsew
rlabel metal1 s 19086 474 19122 815 4 vdd
port 539 nsew
rlabel metal1 s 15822 20224 15858 20565 4 vdd
port 539 nsew
rlabel metal1 s 4110 20224 4146 20565 4 vdd
port 539 nsew
rlabel metal1 s 7854 7875 7890 8216 4 vdd
port 539 nsew
rlabel metal1 s 20814 16565 20850 16906 4 vdd
port 539 nsew
rlabel metal1 s 9582 4424 9618 4765 4 vdd
port 539 nsew
rlabel metal1 s 4590 19434 4626 19775 4 vdd
port 539 nsew
rlabel metal1 s 18318 18935 18354 19276 4 vdd
port 539 nsew
rlabel metal1 s 10350 10744 10386 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 20224 14610 20565 4 vdd
port 539 nsew
rlabel metal1 s 4590 11534 4626 11875 4 vdd
port 539 nsew
rlabel metal1 s 11598 19434 11634 19775 4 vdd
port 539 nsew
rlabel metal1 s 17070 11825 17106 12166 4 vdd
port 539 nsew
rlabel metal1 s 11598 2054 11634 2395 4 vdd
port 539 nsew
rlabel metal1 s 2094 6794 2130 7135 4 vdd
port 539 nsew
rlabel metal1 s 4110 3634 4146 3975 4 vdd
port 539 nsew
rlabel metal1 s 19566 4715 19602 5056 4 vdd
port 539 nsew
rlabel metal1 s 18318 17355 18354 17696 4 vdd
port 539 nsew
rlabel metal1 s 14094 11825 14130 12166 4 vdd
port 539 nsew
rlabel metal1 s 12078 22095 12114 22436 4 vdd
port 539 nsew
rlabel metal1 s 11598 21804 11634 22145 4 vdd
port 539 nsew
rlabel metal1 s 1614 1555 1650 1896 4 vdd
port 539 nsew
rlabel metal1 s 5838 15484 5874 15825 4 vdd
port 539 nsew
rlabel metal1 s 2862 13904 2898 14245 4 vdd
port 539 nsew
rlabel metal1 s 7086 3135 7122 3476 4 vdd
port 539 nsew
rlabel metal1 s 7086 20515 7122 20856 4 vdd
port 539 nsew
rlabel metal1 s 13326 15484 13362 15825 4 vdd
port 539 nsew
rlabel metal1 s 14574 24465 14610 24806 4 vdd
port 539 nsew
rlabel metal1 s 8334 16274 8370 16615 4 vdd
port 539 nsew
rlabel metal1 s 15342 22885 15378 23226 4 vdd
port 539 nsew
rlabel metal1 s 2094 21804 2130 22145 4 vdd
port 539 nsew
rlabel metal1 s 16590 23384 16626 23725 4 vdd
port 539 nsew
rlabel metal1 s 7854 15775 7890 16116 4 vdd
port 539 nsew
rlabel metal1 s 17070 -25 17106 316 4 vdd
port 539 nsew
rlabel metal1 s 10350 5214 10386 5555 4 vdd
port 539 nsew
rlabel metal1 s 6606 22594 6642 22935 4 vdd
port 539 nsew
rlabel metal1 s 20814 5505 20850 5846 4 vdd
port 539 nsew
rlabel metal1 s 10350 14195 10386 14536 4 vdd
port 539 nsew
rlabel metal1 s 15342 3925 15378 4266 4 vdd
port 539 nsew
rlabel metal1 s 14094 17355 14130 17696 4 vdd
port 539 nsew
rlabel metal1 s 6606 4715 6642 5056 4 vdd
port 539 nsew
rlabel metal1 s 1614 12324 1650 12665 4 vdd
port 539 nsew
rlabel metal1 s 20334 6295 20370 6636 4 vdd
port 539 nsew
rlabel metal1 s 10830 7085 10866 7426 4 vdd
port 539 nsew
rlabel metal1 s 12846 9164 12882 9505 4 vdd
port 539 nsew
rlabel metal1 s 4110 19725 4146 20066 4 vdd
port 539 nsew
rlabel metal1 s 5838 18644 5874 18985 4 vdd
port 539 nsew
rlabel metal1 s 9582 10744 9618 11085 4 vdd
port 539 nsew
rlabel metal1 s 1614 22885 1650 23226 4 vdd
port 539 nsew
rlabel metal1 s 20814 1264 20850 1605 4 vdd
port 539 nsew
rlabel metal1 s 1614 765 1650 1106 4 vdd
port 539 nsew
rlabel metal1 s 4590 24465 4626 24806 4 vdd
port 539 nsew
rlabel metal1 s 16590 24465 16626 24806 4 vdd
port 539 nsew
rlabel metal1 s 16590 17355 16626 17696 4 vdd
port 539 nsew
rlabel metal1 s 17070 13405 17106 13746 4 vdd
port 539 nsew
rlabel metal1 s 11598 23384 11634 23725 4 vdd
port 539 nsew
rlabel metal1 s 4590 2345 4626 2686 4 vdd
port 539 nsew
rlabel metal1 s 5358 22885 5394 23226 4 vdd
port 539 nsew
rlabel metal1 s 16590 15775 16626 16116 4 vdd
port 539 nsew
rlabel metal1 s 366 11534 402 11875 4 vdd
port 539 nsew
rlabel metal1 s 9102 18644 9138 18985 4 vdd
port 539 nsew
rlabel metal1 s 5838 765 5874 1106 4 vdd
port 539 nsew
rlabel metal1 s 17838 21014 17874 21355 4 vdd
port 539 nsew
rlabel metal1 s 366 14195 402 14536 4 vdd
port 539 nsew
rlabel metal1 s 4590 13904 4626 14245 4 vdd
port 539 nsew
rlabel metal1 s 17838 7875 17874 8216 4 vdd
port 539 nsew
rlabel metal1 s 19566 24465 19602 24806 4 vdd
port 539 nsew
rlabel metal1 s 6606 9455 6642 9796 4 vdd
port 539 nsew
rlabel metal1 s 2094 4715 2130 5056 4 vdd
port 539 nsew
rlabel metal1 s 3342 1555 3378 1896 4 vdd
port 539 nsew
rlabel metal1 s 12846 13904 12882 14245 4 vdd
port 539 nsew
rlabel metal1 s 15342 3634 15378 3975 4 vdd
port 539 nsew
rlabel metal1 s 846 7584 882 7925 4 vdd
port 539 nsew
rlabel metal1 s 4590 18644 4626 18985 4 vdd
port 539 nsew
rlabel metal1 s 11598 18145 11634 18486 4 vdd
port 539 nsew
rlabel metal1 s 13326 7584 13362 7925 4 vdd
port 539 nsew
rlabel metal1 s 1614 24964 1650 25305 4 vdd
port 539 nsew
rlabel metal1 s 16590 8374 16626 8715 4 vdd
port 539 nsew
rlabel metal1 s 2862 19725 2898 20066 4 vdd
port 539 nsew
rlabel metal1 s 17838 2345 17874 2686 4 vdd
port 539 nsew
rlabel metal1 s 11598 9954 11634 10295 4 vdd
port 539 nsew
rlabel metal1 s 15822 9455 15858 9796 4 vdd
port 539 nsew
rlabel metal1 s 9582 11825 9618 12166 4 vdd
port 539 nsew
rlabel metal1 s 20814 6004 20850 6345 4 vdd
port 539 nsew
rlabel metal1 s 18318 16274 18354 16615 4 vdd
port 539 nsew
rlabel metal1 s 14094 2844 14130 3185 4 vdd
port 539 nsew
rlabel metal1 s 366 22594 402 22935 4 vdd
port 539 nsew
rlabel metal1 s 846 13904 882 14245 4 vdd
port 539 nsew
rlabel metal1 s 17838 6004 17874 6345 4 vdd
port 539 nsew
rlabel metal1 s 11598 10744 11634 11085 4 vdd
port 539 nsew
rlabel metal1 s 19566 21804 19602 22145 4 vdd
port 539 nsew
rlabel metal1 s 7086 17854 7122 18195 4 vdd
port 539 nsew
rlabel metal1 s 15822 12615 15858 12956 4 vdd
port 539 nsew
rlabel metal1 s 19086 20224 19122 20565 4 vdd
port 539 nsew
rlabel metal1 s 9582 6295 9618 6636 4 vdd
port 539 nsew
rlabel metal1 s 16590 12615 16626 12956 4 vdd
port 539 nsew
rlabel metal1 s 846 25255 882 25596 4 vdd
port 539 nsew
rlabel metal1 s 2862 21305 2898 21646 4 vdd
port 539 nsew
rlabel metal1 s 9582 13114 9618 13455 4 vdd
port 539 nsew
rlabel metal1 s 16590 24174 16626 24515 4 vdd
port 539 nsew
rlabel metal1 s 2862 12324 2898 12665 4 vdd
port 539 nsew
rlabel metal1 s 11598 24964 11634 25305 4 vdd
port 539 nsew
rlabel metal1 s 17070 17064 17106 17405 4 vdd
port 539 nsew
rlabel metal1 s 7854 25754 7890 26095 4 vdd
port 539 nsew
rlabel metal1 s 7086 10744 7122 11085 4 vdd
port 539 nsew
rlabel metal1 s 846 24964 882 25305 4 vdd
port 539 nsew
rlabel metal1 s 1614 16565 1650 16906 4 vdd
port 539 nsew
rlabel metal1 s 15342 14694 15378 15035 4 vdd
port 539 nsew
rlabel metal1 s 15342 7584 15378 7925 4 vdd
port 539 nsew
rlabel metal1 s 10350 23384 10386 23725 4 vdd
port 539 nsew
rlabel metal1 s 15822 21804 15858 22145 4 vdd
port 539 nsew
rlabel metal1 s 5358 3925 5394 4266 4 vdd
port 539 nsew
rlabel metal1 s 5358 21305 5394 21646 4 vdd
port 539 nsew
rlabel metal1 s 16590 11534 16626 11875 4 vdd
port 539 nsew
rlabel metal1 s 7086 2345 7122 2686 4 vdd
port 539 nsew
rlabel metal1 s 7086 22095 7122 22436 4 vdd
port 539 nsew
rlabel metal1 s 19086 11534 19122 11875 4 vdd
port 539 nsew
rlabel metal1 s 18318 19434 18354 19775 4 vdd
port 539 nsew
rlabel metal1 s 10830 15484 10866 15825 4 vdd
port 539 nsew
rlabel metal1 s 14574 15775 14610 16116 4 vdd
port 539 nsew
rlabel metal1 s 9582 3634 9618 3975 4 vdd
port 539 nsew
rlabel metal1 s 10350 5505 10386 5846 4 vdd
port 539 nsew
rlabel metal1 s 12078 17064 12114 17405 4 vdd
port 539 nsew
rlabel metal1 s 4590 9164 4626 9505 4 vdd
port 539 nsew
rlabel metal1 s 10350 22594 10386 22935 4 vdd
port 539 nsew
rlabel metal1 s 5358 12615 5394 12956 4 vdd
port 539 nsew
rlabel metal1 s 19566 9954 19602 10295 4 vdd
port 539 nsew
rlabel metal1 s 1614 22095 1650 22436 4 vdd
port 539 nsew
rlabel metal1 s 3342 22885 3378 23226 4 vdd
port 539 nsew
rlabel metal1 s 5358 9954 5394 10295 4 vdd
port 539 nsew
rlabel metal1 s 14094 10744 14130 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 16565 14610 16906 4 vdd
port 539 nsew
rlabel metal1 s 5838 4424 5874 4765 4 vdd
port 539 nsew
rlabel metal1 s 20334 17854 20370 18195 4 vdd
port 539 nsew
rlabel metal1 s 3342 9164 3378 9505 4 vdd
port 539 nsew
rlabel metal1 s 13326 12324 13362 12665 4 vdd
port 539 nsew
rlabel metal1 s 4110 1264 4146 1605 4 vdd
port 539 nsew
rlabel metal1 s 11598 6794 11634 7135 4 vdd
port 539 nsew
rlabel metal1 s 10350 16565 10386 16906 4 vdd
port 539 nsew
rlabel metal1 s 4590 22594 4626 22935 4 vdd
port 539 nsew
rlabel metal1 s 9102 1555 9138 1896 4 vdd
port 539 nsew
rlabel metal1 s 4590 5214 4626 5555 4 vdd
port 539 nsew
rlabel metal1 s 10830 21804 10866 22145 4 vdd
port 539 nsew
rlabel metal1 s 6606 25754 6642 26095 4 vdd
port 539 nsew
rlabel metal1 s 19086 19434 19122 19775 4 vdd
port 539 nsew
rlabel metal1 s 4590 17064 4626 17405 4 vdd
port 539 nsew
rlabel metal1 s 10830 13904 10866 14245 4 vdd
port 539 nsew
rlabel metal1 s 10350 9164 10386 9505 4 vdd
port 539 nsew
rlabel metal1 s 2094 474 2130 815 4 vdd
port 539 nsew
rlabel metal1 s 11598 22885 11634 23226 4 vdd
port 539 nsew
rlabel metal1 s 6606 23384 6642 23725 4 vdd
port 539 nsew
rlabel metal1 s 10350 14694 10386 15035 4 vdd
port 539 nsew
rlabel metal1 s 10830 18644 10866 18985 4 vdd
port 539 nsew
rlabel metal1 s 15342 4424 15378 4765 4 vdd
port 539 nsew
rlabel metal1 s 20334 474 20370 815 4 vdd
port 539 nsew
rlabel metal1 s 5838 13904 5874 14245 4 vdd
port 539 nsew
rlabel metal1 s 9102 3634 9138 3975 4 vdd
port 539 nsew
rlabel metal1 s 14094 765 14130 1106 4 vdd
port 539 nsew
rlabel metal1 s 5838 25255 5874 25596 4 vdd
port 539 nsew
rlabel metal1 s 4590 6295 4626 6636 4 vdd
port 539 nsew
rlabel metal1 s 20814 24465 20850 24806 4 vdd
port 539 nsew
rlabel metal1 s 13326 13904 13362 14245 4 vdd
port 539 nsew
rlabel metal1 s 16590 14985 16626 15326 4 vdd
port 539 nsew
rlabel metal1 s 12078 25255 12114 25596 4 vdd
port 539 nsew
rlabel metal1 s 17838 6794 17874 7135 4 vdd
port 539 nsew
rlabel metal1 s 15342 10744 15378 11085 4 vdd
port 539 nsew
rlabel metal1 s 17838 10245 17874 10586 4 vdd
port 539 nsew
rlabel metal1 s 366 12615 402 12956 4 vdd
port 539 nsew
rlabel metal1 s 366 23675 402 24016 4 vdd
port 539 nsew
rlabel metal1 s 5838 7584 5874 7925 4 vdd
port 539 nsew
rlabel metal1 s 7854 17355 7890 17696 4 vdd
port 539 nsew
rlabel metal1 s 3342 21014 3378 21355 4 vdd
port 539 nsew
rlabel metal1 s 20334 21014 20370 21355 4 vdd
port 539 nsew
rlabel metal1 s 5838 9455 5874 9796 4 vdd
port 539 nsew
rlabel metal1 s 9102 7875 9138 8216 4 vdd
port 539 nsew
rlabel metal1 s 19086 17064 19122 17405 4 vdd
port 539 nsew
rlabel metal1 s 19566 17064 19602 17405 4 vdd
port 539 nsew
rlabel metal1 s 14574 14694 14610 15035 4 vdd
port 539 nsew
rlabel metal1 s 14094 1264 14130 1605 4 vdd
port 539 nsew
rlabel metal1 s 13326 9164 13362 9505 4 vdd
port 539 nsew
rlabel metal1 s 16590 18935 16626 19276 4 vdd
port 539 nsew
rlabel metal1 s 1614 2054 1650 2395 4 vdd
port 539 nsew
rlabel metal1 s 17070 3925 17106 4266 4 vdd
port 539 nsew
rlabel metal1 s 12078 9954 12114 10295 4 vdd
port 539 nsew
rlabel metal1 s 1614 25255 1650 25596 4 vdd
port 539 nsew
rlabel metal1 s 846 10744 882 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 22594 14610 22935 4 vdd
port 539 nsew
rlabel metal1 s 8334 18935 8370 19276 4 vdd
port 539 nsew
rlabel metal1 s 12846 17854 12882 18195 4 vdd
port 539 nsew
rlabel metal1 s 4110 20515 4146 20856 4 vdd
port 539 nsew
rlabel metal1 s 15342 14985 15378 15326 4 vdd
port 539 nsew
rlabel metal1 s 19086 -25 19122 316 4 vdd
port 539 nsew
rlabel metal1 s 18318 12324 18354 12665 4 vdd
port 539 nsew
rlabel metal1 s 7086 11825 7122 12166 4 vdd
port 539 nsew
rlabel metal1 s 11598 9164 11634 9505 4 vdd
port 539 nsew
rlabel metal1 s 20814 18644 20850 18985 4 vdd
port 539 nsew
rlabel metal1 s 7854 7584 7890 7925 4 vdd
port 539 nsew
rlabel metal1 s 12078 8374 12114 8715 4 vdd
port 539 nsew
rlabel metal1 s 15342 8374 15378 8715 4 vdd
port 539 nsew
rlabel metal1 s 7086 7085 7122 7426 4 vdd
port 539 nsew
rlabel metal1 s 13326 474 13362 815 4 vdd
port 539 nsew
rlabel metal1 s 9582 5214 9618 5555 4 vdd
port 539 nsew
rlabel metal1 s 15822 9164 15858 9505 4 vdd
port 539 nsew
rlabel metal1 s 3342 21305 3378 21646 4 vdd
port 539 nsew
rlabel metal1 s 6606 7875 6642 8216 4 vdd
port 539 nsew
rlabel metal1 s 5358 7085 5394 7426 4 vdd
port 539 nsew
rlabel metal1 s 20334 23675 20370 24016 4 vdd
port 539 nsew
rlabel metal1 s 10830 2844 10866 3185 4 vdd
port 539 nsew
rlabel metal1 s 14094 24964 14130 25305 4 vdd
port 539 nsew
rlabel metal1 s 7086 4424 7122 4765 4 vdd
port 539 nsew
rlabel metal1 s 9582 11035 9618 11376 4 vdd
port 539 nsew
rlabel metal1 s 13326 8374 13362 8715 4 vdd
port 539 nsew
rlabel metal1 s 1614 20515 1650 20856 4 vdd
port 539 nsew
rlabel metal1 s 14094 9455 14130 9796 4 vdd
port 539 nsew
rlabel metal1 s 18318 6295 18354 6636 4 vdd
port 539 nsew
rlabel metal1 s 14574 3634 14610 3975 4 vdd
port 539 nsew
rlabel metal1 s 8334 21014 8370 21355 4 vdd
port 539 nsew
rlabel metal1 s 366 21014 402 21355 4 vdd
port 539 nsew
rlabel metal1 s 14574 8665 14610 9006 4 vdd
port 539 nsew
rlabel metal1 s 20334 19434 20370 19775 4 vdd
port 539 nsew
rlabel metal1 s 19566 2844 19602 3185 4 vdd
port 539 nsew
rlabel metal1 s 14574 13114 14610 13455 4 vdd
port 539 nsew
rlabel metal1 s 20814 11534 20850 11875 4 vdd
port 539 nsew
rlabel metal1 s 19086 7584 19122 7925 4 vdd
port 539 nsew
rlabel metal1 s 20334 5505 20370 5846 4 vdd
port 539 nsew
rlabel metal1 s 846 11035 882 11376 4 vdd
port 539 nsew
rlabel metal1 s 14094 18145 14130 18486 4 vdd
port 539 nsew
rlabel metal1 s 20334 11035 20370 11376 4 vdd
port 539 nsew
rlabel metal1 s 18318 13405 18354 13746 4 vdd
port 539 nsew
rlabel metal1 s 846 13114 882 13455 4 vdd
port 539 nsew
rlabel metal1 s 10830 4424 10866 4765 4 vdd
port 539 nsew
rlabel metal1 s 2094 16565 2130 16906 4 vdd
port 539 nsew
rlabel metal1 s 5838 17064 5874 17405 4 vdd
port 539 nsew
rlabel metal1 s 2862 20515 2898 20856 4 vdd
port 539 nsew
rlabel metal1 s 17070 765 17106 1106 4 vdd
port 539 nsew
rlabel metal1 s 19566 5214 19602 5555 4 vdd
port 539 nsew
rlabel metal1 s 16590 17854 16626 18195 4 vdd
port 539 nsew
rlabel metal1 s 10350 6295 10386 6636 4 vdd
port 539 nsew
rlabel metal1 s 2862 -25 2898 316 4 vdd
port 539 nsew
rlabel metal1 s 3342 11035 3378 11376 4 vdd
port 539 nsew
rlabel metal1 s 10830 -25 10866 316 4 vdd
port 539 nsew
rlabel metal1 s 19566 24964 19602 25305 4 vdd
port 539 nsew
rlabel metal1 s 17070 21014 17106 21355 4 vdd
port 539 nsew
rlabel metal1 s 13326 5505 13362 5846 4 vdd
port 539 nsew
rlabel metal1 s 17070 16274 17106 16615 4 vdd
port 539 nsew
rlabel metal1 s 16590 9954 16626 10295 4 vdd
port 539 nsew
rlabel metal1 s 2094 12324 2130 12665 4 vdd
port 539 nsew
rlabel metal1 s 15342 9455 15378 9796 4 vdd
port 539 nsew
rlabel metal1 s 7086 23675 7122 24016 4 vdd
port 539 nsew
rlabel metal1 s 17070 16565 17106 16906 4 vdd
port 539 nsew
rlabel metal1 s 6606 10245 6642 10586 4 vdd
port 539 nsew
rlabel metal1 s 9582 765 9618 1106 4 vdd
port 539 nsew
rlabel metal1 s 20334 25255 20370 25596 4 vdd
port 539 nsew
rlabel metal1 s 5838 20224 5874 20565 4 vdd
port 539 nsew
rlabel metal1 s 2862 24465 2898 24806 4 vdd
port 539 nsew
rlabel metal1 s 11598 765 11634 1106 4 vdd
port 539 nsew
rlabel metal1 s 10830 22885 10866 23226 4 vdd
port 539 nsew
rlabel metal1 s 7086 18145 7122 18486 4 vdd
port 539 nsew
rlabel metal1 s 14094 6794 14130 7135 4 vdd
port 539 nsew
rlabel metal1 s 15822 14985 15858 15326 4 vdd
port 539 nsew
rlabel metal1 s 11598 3925 11634 4266 4 vdd
port 539 nsew
rlabel metal1 s 17070 5214 17106 5555 4 vdd
port 539 nsew
rlabel metal1 s 4590 765 4626 1106 4 vdd
port 539 nsew
rlabel metal1 s 13326 7875 13362 8216 4 vdd
port 539 nsew
rlabel metal1 s 2862 7875 2898 8216 4 vdd
port 539 nsew
rlabel metal1 s 16590 22095 16626 22436 4 vdd
port 539 nsew
rlabel metal1 s 16590 1264 16626 1605 4 vdd
port 539 nsew
rlabel metal1 s 12078 24964 12114 25305 4 vdd
port 539 nsew
rlabel metal1 s 19086 3135 19122 3476 4 vdd
port 539 nsew
rlabel metal1 s 8334 20224 8370 20565 4 vdd
port 539 nsew
rlabel metal1 s 14574 19434 14610 19775 4 vdd
port 539 nsew
rlabel metal1 s 19566 2054 19602 2395 4 vdd
port 539 nsew
rlabel metal1 s 366 15484 402 15825 4 vdd
port 539 nsew
rlabel metal1 s 7086 12615 7122 12956 4 vdd
port 539 nsew
rlabel metal1 s 16590 22594 16626 22935 4 vdd
port 539 nsew
rlabel metal1 s 14094 21804 14130 22145 4 vdd
port 539 nsew
rlabel metal1 s 10350 10245 10386 10586 4 vdd
port 539 nsew
rlabel metal1 s 12078 24174 12114 24515 4 vdd
port 539 nsew
rlabel metal1 s 9582 11534 9618 11875 4 vdd
port 539 nsew
rlabel metal1 s 10350 7085 10386 7426 4 vdd
port 539 nsew
rlabel metal1 s 2094 11534 2130 11875 4 vdd
port 539 nsew
rlabel metal1 s 2862 15775 2898 16116 4 vdd
port 539 nsew
rlabel metal1 s 6606 3135 6642 3476 4 vdd
port 539 nsew
rlabel metal1 s 17070 18145 17106 18486 4 vdd
port 539 nsew
rlabel metal1 s 15342 13114 15378 13455 4 vdd
port 539 nsew
rlabel metal1 s 7086 3634 7122 3975 4 vdd
port 539 nsew
rlabel metal1 s 19086 23675 19122 24016 4 vdd
port 539 nsew
rlabel metal1 s 7854 5505 7890 5846 4 vdd
port 539 nsew
rlabel metal1 s 18318 9954 18354 10295 4 vdd
port 539 nsew
rlabel metal1 s 366 3925 402 4266 4 vdd
port 539 nsew
rlabel metal1 s 10350 -25 10386 316 4 vdd
port 539 nsew
rlabel metal1 s 19086 21305 19122 21646 4 vdd
port 539 nsew
rlabel metal1 s 17070 3634 17106 3975 4 vdd
port 539 nsew
rlabel metal1 s 17070 7875 17106 8216 4 vdd
port 539 nsew
rlabel metal1 s 1614 2844 1650 3185 4 vdd
port 539 nsew
rlabel metal1 s 17838 24964 17874 25305 4 vdd
port 539 nsew
rlabel metal1 s 5838 2345 5874 2686 4 vdd
port 539 nsew
rlabel metal1 s 12078 11825 12114 12166 4 vdd
port 539 nsew
rlabel metal1 s 14574 7085 14610 7426 4 vdd
port 539 nsew
rlabel metal1 s 5838 23384 5874 23725 4 vdd
port 539 nsew
rlabel metal1 s 11598 15484 11634 15825 4 vdd
port 539 nsew
rlabel metal1 s 846 1264 882 1605 4 vdd
port 539 nsew
rlabel metal1 s 846 12615 882 12956 4 vdd
port 539 nsew
rlabel metal1 s 15822 22885 15858 23226 4 vdd
port 539 nsew
rlabel metal1 s 7086 14985 7122 15326 4 vdd
port 539 nsew
rlabel metal1 s 9102 24174 9138 24515 4 vdd
port 539 nsew
rlabel metal1 s 9582 3925 9618 4266 4 vdd
port 539 nsew
rlabel metal1 s 5838 24465 5874 24806 4 vdd
port 539 nsew
rlabel metal1 s 12846 10245 12882 10586 4 vdd
port 539 nsew
rlabel metal1 s 1614 13405 1650 13746 4 vdd
port 539 nsew
rlabel metal1 s 12846 16274 12882 16615 4 vdd
port 539 nsew
rlabel metal1 s 6606 17355 6642 17696 4 vdd
port 539 nsew
rlabel metal1 s 20334 10744 20370 11085 4 vdd
port 539 nsew
rlabel metal1 s 366 1555 402 1896 4 vdd
port 539 nsew
rlabel metal1 s 12078 5214 12114 5555 4 vdd
port 539 nsew
rlabel metal1 s 15822 19434 15858 19775 4 vdd
port 539 nsew
rlabel metal1 s 4110 24465 4146 24806 4 vdd
port 539 nsew
rlabel metal1 s 18318 1264 18354 1605 4 vdd
port 539 nsew
rlabel metal1 s 7086 4715 7122 5056 4 vdd
port 539 nsew
rlabel metal1 s 13326 9455 13362 9796 4 vdd
port 539 nsew
rlabel metal1 s 9102 3135 9138 3476 4 vdd
port 539 nsew
rlabel metal1 s 17070 3135 17106 3476 4 vdd
port 539 nsew
rlabel metal1 s 2862 13114 2898 13455 4 vdd
port 539 nsew
rlabel metal1 s 19566 1555 19602 1896 4 vdd
port 539 nsew
rlabel metal1 s 3342 4715 3378 5056 4 vdd
port 539 nsew
rlabel metal1 s 19086 11825 19122 12166 4 vdd
port 539 nsew
rlabel metal1 s 4110 7085 4146 7426 4 vdd
port 539 nsew
rlabel metal1 s 3342 14195 3378 14536 4 vdd
port 539 nsew
rlabel metal1 s 13326 17854 13362 18195 4 vdd
port 539 nsew
rlabel metal1 s 13326 13405 13362 13746 4 vdd
port 539 nsew
rlabel metal1 s 14574 6794 14610 7135 4 vdd
port 539 nsew
rlabel metal1 s 5838 21014 5874 21355 4 vdd
port 539 nsew
rlabel metal1 s 19566 22594 19602 22935 4 vdd
port 539 nsew
rlabel metal1 s 14574 6295 14610 6636 4 vdd
port 539 nsew
rlabel metal1 s 2094 11825 2130 12166 4 vdd
port 539 nsew
rlabel metal1 s 846 5505 882 5846 4 vdd
port 539 nsew
rlabel metal1 s 12846 19434 12882 19775 4 vdd
port 539 nsew
rlabel metal1 s 19566 7584 19602 7925 4 vdd
port 539 nsew
rlabel metal1 s 14094 3925 14130 4266 4 vdd
port 539 nsew
rlabel metal1 s 16590 9455 16626 9796 4 vdd
port 539 nsew
rlabel metal1 s 9102 6794 9138 7135 4 vdd
port 539 nsew
rlabel metal1 s 9582 22885 9618 23226 4 vdd
port 539 nsew
rlabel metal1 s 7086 24964 7122 25305 4 vdd
port 539 nsew
rlabel metal1 s 20334 6794 20370 7135 4 vdd
port 539 nsew
rlabel metal1 s 20814 21305 20850 21646 4 vdd
port 539 nsew
rlabel metal1 s 5838 11825 5874 12166 4 vdd
port 539 nsew
rlabel metal1 s 19566 20515 19602 20856 4 vdd
port 539 nsew
rlabel metal1 s 20814 14694 20850 15035 4 vdd
port 539 nsew
rlabel metal1 s 12846 25754 12882 26095 4 vdd
port 539 nsew
rlabel metal1 s 5358 12324 5394 12665 4 vdd
port 539 nsew
rlabel metal1 s 4590 22095 4626 22436 4 vdd
port 539 nsew
rlabel metal1 s 1614 17064 1650 17405 4 vdd
port 539 nsew
rlabel metal1 s 7854 14694 7890 15035 4 vdd
port 539 nsew
rlabel metal1 s 9102 13114 9138 13455 4 vdd
port 539 nsew
rlabel metal1 s 5838 11035 5874 11376 4 vdd
port 539 nsew
rlabel metal1 s 5358 5214 5394 5555 4 vdd
port 539 nsew
rlabel metal1 s 9102 15484 9138 15825 4 vdd
port 539 nsew
rlabel metal1 s 1614 9954 1650 10295 4 vdd
port 539 nsew
rlabel metal1 s 7086 14694 7122 15035 4 vdd
port 539 nsew
rlabel metal1 s 6606 11825 6642 12166 4 vdd
port 539 nsew
rlabel metal1 s 8334 24174 8370 24515 4 vdd
port 539 nsew
rlabel metal1 s 11598 11534 11634 11875 4 vdd
port 539 nsew
rlabel metal1 s 5838 19434 5874 19775 4 vdd
port 539 nsew
rlabel metal1 s 19086 13405 19122 13746 4 vdd
port 539 nsew
rlabel metal1 s 10350 18145 10386 18486 4 vdd
port 539 nsew
rlabel metal1 s 11598 4715 11634 5056 4 vdd
port 539 nsew
rlabel metal1 s 14094 14195 14130 14536 4 vdd
port 539 nsew
rlabel metal1 s 10350 18644 10386 18985 4 vdd
port 539 nsew
rlabel metal1 s 12078 3925 12114 4266 4 vdd
port 539 nsew
rlabel metal1 s 12078 2844 12114 3185 4 vdd
port 539 nsew
rlabel metal1 s 17838 13114 17874 13455 4 vdd
port 539 nsew
rlabel metal1 s 1614 1264 1650 1605 4 vdd
port 539 nsew
rlabel metal1 s 7854 16274 7890 16615 4 vdd
port 539 nsew
rlabel metal1 s 13326 16565 13362 16906 4 vdd
port 539 nsew
rlabel metal1 s 9582 474 9618 815 4 vdd
port 539 nsew
rlabel metal1 s 15822 15775 15858 16116 4 vdd
port 539 nsew
rlabel metal1 s 16590 7875 16626 8216 4 vdd
port 539 nsew
rlabel metal1 s 2862 2054 2898 2395 4 vdd
port 539 nsew
rlabel metal1 s 10350 6004 10386 6345 4 vdd
port 539 nsew
rlabel metal1 s 366 17854 402 18195 4 vdd
port 539 nsew
rlabel metal1 s 14574 15484 14610 15825 4 vdd
port 539 nsew
rlabel metal1 s 7854 13405 7890 13746 4 vdd
port 539 nsew
rlabel metal1 s 8334 474 8370 815 4 vdd
port 539 nsew
rlabel metal1 s 9102 21305 9138 21646 4 vdd
port 539 nsew
rlabel metal1 s 2094 13405 2130 13746 4 vdd
port 539 nsew
rlabel metal1 s 4590 18145 4626 18486 4 vdd
port 539 nsew
rlabel metal1 s 2094 3135 2130 3476 4 vdd
port 539 nsew
rlabel metal1 s 3342 10744 3378 11085 4 vdd
port 539 nsew
rlabel metal1 s 20334 2054 20370 2395 4 vdd
port 539 nsew
rlabel metal1 s 16590 24964 16626 25305 4 vdd
port 539 nsew
rlabel metal1 s 18318 21305 18354 21646 4 vdd
port 539 nsew
rlabel metal1 s 4110 9164 4146 9505 4 vdd
port 539 nsew
rlabel metal1 s 13326 21804 13362 22145 4 vdd
port 539 nsew
rlabel metal1 s 9102 22095 9138 22436 4 vdd
port 539 nsew
rlabel metal1 s 2862 11534 2898 11875 4 vdd
port 539 nsew
rlabel metal1 s 5838 8374 5874 8715 4 vdd
port 539 nsew
rlabel metal1 s 12846 15484 12882 15825 4 vdd
port 539 nsew
rlabel metal1 s 7854 13114 7890 13455 4 vdd
port 539 nsew
rlabel metal1 s 366 765 402 1106 4 vdd
port 539 nsew
rlabel metal1 s 15342 21014 15378 21355 4 vdd
port 539 nsew
rlabel metal1 s 3342 2054 3378 2395 4 vdd
port 539 nsew
rlabel metal1 s 8334 14195 8370 14536 4 vdd
port 539 nsew
rlabel metal1 s 7086 11534 7122 11875 4 vdd
port 539 nsew
rlabel metal1 s 6606 6794 6642 7135 4 vdd
port 539 nsew
rlabel metal1 s 2862 5505 2898 5846 4 vdd
port 539 nsew
rlabel metal1 s 15342 17854 15378 18195 4 vdd
port 539 nsew
rlabel metal1 s 16590 10744 16626 11085 4 vdd
port 539 nsew
rlabel metal1 s 18318 3135 18354 3476 4 vdd
port 539 nsew
rlabel metal1 s 5838 10744 5874 11085 4 vdd
port 539 nsew
rlabel metal1 s 14094 9954 14130 10295 4 vdd
port 539 nsew
rlabel metal1 s 9582 14694 9618 15035 4 vdd
port 539 nsew
rlabel metal1 s 13326 2844 13362 3185 4 vdd
port 539 nsew
rlabel metal1 s 1614 21804 1650 22145 4 vdd
port 539 nsew
rlabel metal1 s 7854 14195 7890 14536 4 vdd
port 539 nsew
rlabel metal1 s 20334 8374 20370 8715 4 vdd
port 539 nsew
rlabel metal1 s 2094 9954 2130 10295 4 vdd
port 539 nsew
rlabel metal1 s 2094 2844 2130 3185 4 vdd
port 539 nsew
rlabel metal1 s 16590 23675 16626 24016 4 vdd
port 539 nsew
rlabel metal1 s 20814 15775 20850 16116 4 vdd
port 539 nsew
rlabel metal1 s 14094 15775 14130 16116 4 vdd
port 539 nsew
rlabel metal1 s 11598 10245 11634 10586 4 vdd
port 539 nsew
rlabel metal1 s 20334 24964 20370 25305 4 vdd
port 539 nsew
rlabel metal1 s 2862 21014 2898 21355 4 vdd
port 539 nsew
rlabel metal1 s 19566 20224 19602 20565 4 vdd
port 539 nsew
rlabel metal1 s 10350 9954 10386 10295 4 vdd
port 539 nsew
rlabel metal1 s 15342 1555 15378 1896 4 vdd
port 539 nsew
rlabel metal1 s 12846 19725 12882 20066 4 vdd
port 539 nsew
rlabel metal1 s 12846 18644 12882 18985 4 vdd
port 539 nsew
rlabel metal1 s 6606 14985 6642 15326 4 vdd
port 539 nsew
rlabel metal1 s 19566 10744 19602 11085 4 vdd
port 539 nsew
rlabel metal1 s 14574 4424 14610 4765 4 vdd
port 539 nsew
rlabel metal1 s 15822 21305 15858 21646 4 vdd
port 539 nsew
rlabel metal1 s 15822 8374 15858 8715 4 vdd
port 539 nsew
rlabel metal1 s 17070 22885 17106 23226 4 vdd
port 539 nsew
rlabel metal1 s 10830 8374 10866 8715 4 vdd
port 539 nsew
rlabel metal1 s 20814 11825 20850 12166 4 vdd
port 539 nsew
rlabel metal1 s 846 18935 882 19276 4 vdd
port 539 nsew
rlabel metal1 s 19566 18935 19602 19276 4 vdd
port 539 nsew
rlabel metal1 s 8334 10245 8370 10586 4 vdd
port 539 nsew
rlabel metal1 s 20814 16274 20850 16615 4 vdd
port 539 nsew
rlabel metal1 s 9582 23384 9618 23725 4 vdd
port 539 nsew
rlabel metal1 s 10350 3135 10386 3476 4 vdd
port 539 nsew
rlabel metal1 s 14574 18935 14610 19276 4 vdd
port 539 nsew
rlabel metal1 s 13326 6794 13362 7135 4 vdd
port 539 nsew
rlabel metal1 s 2094 8374 2130 8715 4 vdd
port 539 nsew
rlabel metal1 s 8334 25255 8370 25596 4 vdd
port 539 nsew
rlabel metal1 s 20814 -25 20850 316 4 vdd
port 539 nsew
rlabel metal1 s 16590 4715 16626 5056 4 vdd
port 539 nsew
rlabel metal1 s 9102 2054 9138 2395 4 vdd
port 539 nsew
rlabel metal1 s 19086 22885 19122 23226 4 vdd
port 539 nsew
rlabel metal1 s 15342 20515 15378 20856 4 vdd
port 539 nsew
rlabel metal1 s 1614 23675 1650 24016 4 vdd
port 539 nsew
rlabel metal1 s 14094 1555 14130 1896 4 vdd
port 539 nsew
rlabel metal1 s 12846 17355 12882 17696 4 vdd
port 539 nsew
rlabel metal1 s 366 22095 402 22436 4 vdd
port 539 nsew
rlabel metal1 s 5838 17355 5874 17696 4 vdd
port 539 nsew
rlabel metal1 s 12846 6004 12882 6345 4 vdd
port 539 nsew
rlabel metal1 s 10830 4715 10866 5056 4 vdd
port 539 nsew
rlabel metal1 s 8334 17064 8370 17405 4 vdd
port 539 nsew
rlabel metal1 s 15822 10744 15858 11085 4 vdd
port 539 nsew
rlabel metal1 s 12078 18935 12114 19276 4 vdd
port 539 nsew
rlabel metal1 s 13326 7085 13362 7426 4 vdd
port 539 nsew
rlabel metal1 s 4590 12324 4626 12665 4 vdd
port 539 nsew
rlabel metal1 s 16590 14694 16626 15035 4 vdd
port 539 nsew
rlabel metal1 s 2862 19434 2898 19775 4 vdd
port 539 nsew
rlabel metal1 s 17838 11825 17874 12166 4 vdd
port 539 nsew
rlabel metal1 s 10350 15775 10386 16116 4 vdd
port 539 nsew
rlabel metal1 s 20334 7875 20370 8216 4 vdd
port 539 nsew
rlabel metal1 s 5838 5214 5874 5555 4 vdd
port 539 nsew
rlabel metal1 s 6606 12324 6642 12665 4 vdd
port 539 nsew
rlabel metal1 s 3342 17854 3378 18195 4 vdd
port 539 nsew
rlabel metal1 s 20334 3925 20370 4266 4 vdd
port 539 nsew
rlabel metal1 s 5358 15775 5394 16116 4 vdd
port 539 nsew
rlabel metal1 s 6606 17064 6642 17405 4 vdd
port 539 nsew
rlabel metal1 s 4110 7875 4146 8216 4 vdd
port 539 nsew
rlabel metal1 s 8334 17854 8370 18195 4 vdd
port 539 nsew
rlabel metal1 s 10830 21305 10866 21646 4 vdd
port 539 nsew
rlabel metal1 s 366 14694 402 15035 4 vdd
port 539 nsew
rlabel metal1 s 15822 23675 15858 24016 4 vdd
port 539 nsew
rlabel metal1 s 14094 16565 14130 16906 4 vdd
port 539 nsew
rlabel metal1 s 9102 14985 9138 15326 4 vdd
port 539 nsew
rlabel metal1 s 846 2054 882 2395 4 vdd
port 539 nsew
rlabel metal1 s 9102 17064 9138 17405 4 vdd
port 539 nsew
rlabel metal1 s 1614 -25 1650 316 4 vdd
port 539 nsew
rlabel metal1 s 15822 17355 15858 17696 4 vdd
port 539 nsew
rlabel metal1 s 20814 7584 20850 7925 4 vdd
port 539 nsew
rlabel metal1 s 19566 17854 19602 18195 4 vdd
port 539 nsew
rlabel metal1 s 2094 25255 2130 25596 4 vdd
port 539 nsew
rlabel metal1 s 1614 17355 1650 17696 4 vdd
port 539 nsew
rlabel metal1 s 6606 6295 6642 6636 4 vdd
port 539 nsew
rlabel metal1 s 15342 12324 15378 12665 4 vdd
port 539 nsew
rlabel metal1 s 17070 23675 17106 24016 4 vdd
port 539 nsew
rlabel metal1 s 7854 12615 7890 12956 4 vdd
port 539 nsew
rlabel metal1 s 8334 19434 8370 19775 4 vdd
port 539 nsew
rlabel metal1 s 6606 16274 6642 16615 4 vdd
port 539 nsew
rlabel metal1 s 19566 16565 19602 16906 4 vdd
port 539 nsew
rlabel metal1 s 9102 2345 9138 2686 4 vdd
port 539 nsew
rlabel metal1 s 7854 7085 7890 7426 4 vdd
port 539 nsew
rlabel metal1 s 9102 11825 9138 12166 4 vdd
port 539 nsew
rlabel metal1 s 15822 2345 15858 2686 4 vdd
port 539 nsew
rlabel metal1 s 846 17854 882 18195 4 vdd
port 539 nsew
rlabel metal1 s 2094 10245 2130 10586 4 vdd
port 539 nsew
rlabel metal1 s 11598 5505 11634 5846 4 vdd
port 539 nsew
rlabel metal1 s 17070 24174 17106 24515 4 vdd
port 539 nsew
rlabel metal1 s 10830 10245 10866 10586 4 vdd
port 539 nsew
rlabel metal1 s 3342 17355 3378 17696 4 vdd
port 539 nsew
rlabel metal1 s 5838 11534 5874 11875 4 vdd
port 539 nsew
rlabel metal1 s 846 6794 882 7135 4 vdd
port 539 nsew
rlabel metal1 s 4110 15775 4146 16116 4 vdd
port 539 nsew
rlabel metal1 s 19566 4424 19602 4765 4 vdd
port 539 nsew
rlabel metal1 s 3342 474 3378 815 4 vdd
port 539 nsew
rlabel metal1 s 2094 -25 2130 316 4 vdd
port 539 nsew
rlabel metal1 s 17838 12324 17874 12665 4 vdd
port 539 nsew
rlabel metal1 s 10830 24174 10866 24515 4 vdd
port 539 nsew
rlabel metal1 s 6606 22885 6642 23226 4 vdd
port 539 nsew
rlabel metal1 s 19086 2844 19122 3185 4 vdd
port 539 nsew
rlabel metal1 s 17838 25255 17874 25596 4 vdd
port 539 nsew
rlabel metal1 s 11598 25255 11634 25596 4 vdd
port 539 nsew
rlabel metal1 s 12078 4715 12114 5056 4 vdd
port 539 nsew
rlabel metal1 s 9102 13904 9138 14245 4 vdd
port 539 nsew
rlabel metal1 s 10830 474 10866 815 4 vdd
port 539 nsew
rlabel metal1 s 9582 20224 9618 20565 4 vdd
port 539 nsew
rlabel metal1 s 12846 3135 12882 3476 4 vdd
port 539 nsew
rlabel metal1 s 13326 17064 13362 17405 4 vdd
port 539 nsew
rlabel metal1 s 13326 2054 13362 2395 4 vdd
port 539 nsew
rlabel metal1 s 4110 7584 4146 7925 4 vdd
port 539 nsew
rlabel metal1 s 15342 25255 15378 25596 4 vdd
port 539 nsew
rlabel metal1 s 13326 11035 13362 11376 4 vdd
port 539 nsew
rlabel metal1 s 366 10245 402 10586 4 vdd
port 539 nsew
rlabel metal1 s 1614 12615 1650 12956 4 vdd
port 539 nsew
rlabel metal1 s 11598 2844 11634 3185 4 vdd
port 539 nsew
rlabel metal1 s 14094 4424 14130 4765 4 vdd
port 539 nsew
rlabel metal1 s 4110 15484 4146 15825 4 vdd
port 539 nsew
rlabel metal1 s 12846 1555 12882 1896 4 vdd
port 539 nsew
rlabel metal1 s 13326 10245 13362 10586 4 vdd
port 539 nsew
rlabel metal1 s 12846 2054 12882 2395 4 vdd
port 539 nsew
rlabel metal1 s 6606 10744 6642 11085 4 vdd
port 539 nsew
rlabel metal1 s 19086 7875 19122 8216 4 vdd
port 539 nsew
rlabel metal1 s 19086 25255 19122 25596 4 vdd
port 539 nsew
rlabel metal1 s 17070 14195 17106 14536 4 vdd
port 539 nsew
rlabel metal1 s 19566 13405 19602 13746 4 vdd
port 539 nsew
rlabel metal1 s 19566 15775 19602 16116 4 vdd
port 539 nsew
rlabel metal1 s 846 3135 882 3476 4 vdd
port 539 nsew
rlabel metal1 s 20814 19725 20850 20066 4 vdd
port 539 nsew
rlabel metal1 s 9582 7875 9618 8216 4 vdd
port 539 nsew
rlabel metal1 s 846 25754 882 26095 4 vdd
port 539 nsew
rlabel metal1 s 19566 7875 19602 8216 4 vdd
port 539 nsew
rlabel metal1 s 366 2054 402 2395 4 vdd
port 539 nsew
rlabel metal1 s 7086 10245 7122 10586 4 vdd
port 539 nsew
rlabel metal1 s 2862 11825 2898 12166 4 vdd
port 539 nsew
rlabel metal1 s 17838 7584 17874 7925 4 vdd
port 539 nsew
rlabel metal1 s 5838 21305 5874 21646 4 vdd
port 539 nsew
rlabel metal1 s 20814 8374 20850 8715 4 vdd
port 539 nsew
rlabel metal1 s 18318 7875 18354 8216 4 vdd
port 539 nsew
rlabel metal1 s 16590 16274 16626 16615 4 vdd
port 539 nsew
rlabel metal1 s 19086 9164 19122 9505 4 vdd
port 539 nsew
rlabel metal1 s 7854 8374 7890 8715 4 vdd
port 539 nsew
rlabel metal1 s 20814 765 20850 1106 4 vdd
port 539 nsew
rlabel metal1 s 17838 21804 17874 22145 4 vdd
port 539 nsew
rlabel metal1 s 9582 1555 9618 1896 4 vdd
port 539 nsew
rlabel metal1 s 7086 18644 7122 18985 4 vdd
port 539 nsew
rlabel metal1 s 14094 13114 14130 13455 4 vdd
port 539 nsew
rlabel metal1 s 15342 11825 15378 12166 4 vdd
port 539 nsew
rlabel metal1 s 366 13405 402 13746 4 vdd
port 539 nsew
rlabel metal1 s 15822 16565 15858 16906 4 vdd
port 539 nsew
rlabel metal1 s 15342 24465 15378 24806 4 vdd
port 539 nsew
rlabel metal1 s 15342 17064 15378 17405 4 vdd
port 539 nsew
rlabel metal1 s 15342 24174 15378 24515 4 vdd
port 539 nsew
rlabel metal1 s 13326 24174 13362 24515 4 vdd
port 539 nsew
rlabel metal1 s 15822 9954 15858 10295 4 vdd
port 539 nsew
rlabel metal1 s 2862 22095 2898 22436 4 vdd
port 539 nsew
rlabel metal1 s 5358 765 5394 1106 4 vdd
port 539 nsew
rlabel metal1 s 8334 13114 8370 13455 4 vdd
port 539 nsew
rlabel metal1 s 4110 5505 4146 5846 4 vdd
port 539 nsew
rlabel metal1 s 366 7584 402 7925 4 vdd
port 539 nsew
rlabel metal1 s 13326 5214 13362 5555 4 vdd
port 539 nsew
rlabel metal1 s 8334 4424 8370 4765 4 vdd
port 539 nsew
rlabel metal1 s 14574 8374 14610 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 4424 9138 4765 4 vdd
port 539 nsew
rlabel metal1 s 12078 17355 12114 17696 4 vdd
port 539 nsew
rlabel metal1 s 7086 7875 7122 8216 4 vdd
port 539 nsew
rlabel metal1 s 10830 19725 10866 20066 4 vdd
port 539 nsew
rlabel metal1 s 19566 -25 19602 316 4 vdd
port 539 nsew
rlabel metal1 s 2862 22594 2898 22935 4 vdd
port 539 nsew
rlabel metal1 s 9102 765 9138 1106 4 vdd
port 539 nsew
rlabel metal1 s 2094 5214 2130 5555 4 vdd
port 539 nsew
rlabel metal1 s 19566 11534 19602 11875 4 vdd
port 539 nsew
rlabel metal1 s 10350 4424 10386 4765 4 vdd
port 539 nsew
rlabel metal1 s 5358 1264 5394 1605 4 vdd
port 539 nsew
rlabel metal1 s 10830 11825 10866 12166 4 vdd
port 539 nsew
rlabel metal1 s 7086 5214 7122 5555 4 vdd
port 539 nsew
rlabel metal1 s 11598 8665 11634 9006 4 vdd
port 539 nsew
rlabel metal1 s 13326 10744 13362 11085 4 vdd
port 539 nsew
rlabel metal1 s 15342 2345 15378 2686 4 vdd
port 539 nsew
rlabel metal1 s 13326 4424 13362 4765 4 vdd
port 539 nsew
rlabel metal1 s 15342 11534 15378 11875 4 vdd
port 539 nsew
rlabel metal1 s 846 16274 882 16615 4 vdd
port 539 nsew
rlabel metal1 s 8334 5505 8370 5846 4 vdd
port 539 nsew
rlabel metal1 s 17838 5505 17874 5846 4 vdd
port 539 nsew
rlabel metal1 s 5838 16565 5874 16906 4 vdd
port 539 nsew
rlabel metal1 s 8334 8665 8370 9006 4 vdd
port 539 nsew
rlabel metal1 s 7854 21014 7890 21355 4 vdd
port 539 nsew
rlabel metal1 s 4110 23675 4146 24016 4 vdd
port 539 nsew
rlabel metal1 s 18318 13904 18354 14245 4 vdd
port 539 nsew
rlabel metal1 s 5358 7875 5394 8216 4 vdd
port 539 nsew
rlabel metal1 s 4590 1264 4626 1605 4 vdd
port 539 nsew
rlabel metal1 s 366 12324 402 12665 4 vdd
port 539 nsew
rlabel metal1 s 5358 6295 5394 6636 4 vdd
port 539 nsew
rlabel metal1 s 5838 10245 5874 10586 4 vdd
port 539 nsew
rlabel metal1 s 4110 23384 4146 23725 4 vdd
port 539 nsew
rlabel metal1 s 15342 19434 15378 19775 4 vdd
port 539 nsew
rlabel metal1 s 10350 3634 10386 3975 4 vdd
port 539 nsew
rlabel metal1 s 12846 7584 12882 7925 4 vdd
port 539 nsew
rlabel metal1 s 1614 15484 1650 15825 4 vdd
port 539 nsew
rlabel metal1 s 20334 11534 20370 11875 4 vdd
port 539 nsew
rlabel metal1 s 8334 12324 8370 12665 4 vdd
port 539 nsew
rlabel metal1 s 9102 6004 9138 6345 4 vdd
port 539 nsew
rlabel metal1 s 3342 6794 3378 7135 4 vdd
port 539 nsew
rlabel metal1 s 4590 13405 4626 13746 4 vdd
port 539 nsew
rlabel metal1 s 13326 22594 13362 22935 4 vdd
port 539 nsew
rlabel metal1 s 5838 22594 5874 22935 4 vdd
port 539 nsew
rlabel metal1 s 366 2345 402 2686 4 vdd
port 539 nsew
rlabel metal1 s 20334 2844 20370 3185 4 vdd
port 539 nsew
rlabel metal1 s 12078 10744 12114 11085 4 vdd
port 539 nsew
rlabel metal1 s 7086 17355 7122 17696 4 vdd
port 539 nsew
rlabel metal1 s 3342 12324 3378 12665 4 vdd
port 539 nsew
rlabel metal1 s 14094 7875 14130 8216 4 vdd
port 539 nsew
rlabel metal1 s 4590 12615 4626 12956 4 vdd
port 539 nsew
rlabel metal1 s 846 765 882 1106 4 vdd
port 539 nsew
rlabel metal1 s 5358 13114 5394 13455 4 vdd
port 539 nsew
rlabel metal1 s 7854 12324 7890 12665 4 vdd
port 539 nsew
rlabel metal1 s 15822 10245 15858 10586 4 vdd
port 539 nsew
rlabel metal1 s 1614 11534 1650 11875 4 vdd
port 539 nsew
rlabel metal1 s 20334 13405 20370 13746 4 vdd
port 539 nsew
rlabel metal1 s 6606 2844 6642 3185 4 vdd
port 539 nsew
rlabel metal1 s 15342 6004 15378 6345 4 vdd
port 539 nsew
rlabel metal1 s 11598 12615 11634 12956 4 vdd
port 539 nsew
rlabel metal1 s 846 18644 882 18985 4 vdd
port 539 nsew
rlabel metal1 s 11598 -25 11634 316 4 vdd
port 539 nsew
rlabel metal1 s 2094 11035 2130 11376 4 vdd
port 539 nsew
rlabel metal1 s 2862 3925 2898 4266 4 vdd
port 539 nsew
rlabel metal1 s 19086 3925 19122 4266 4 vdd
port 539 nsew
rlabel metal1 s 19566 2345 19602 2686 4 vdd
port 539 nsew
rlabel metal1 s 13326 3135 13362 3476 4 vdd
port 539 nsew
rlabel metal1 s 10830 16274 10866 16615 4 vdd
port 539 nsew
rlabel metal1 s 20334 25754 20370 26095 4 vdd
port 539 nsew
rlabel metal1 s 14094 14694 14130 15035 4 vdd
port 539 nsew
rlabel metal1 s 10350 11534 10386 11875 4 vdd
port 539 nsew
rlabel metal1 s 2094 21014 2130 21355 4 vdd
port 539 nsew
rlabel metal1 s 366 1264 402 1605 4 vdd
port 539 nsew
rlabel metal1 s 12078 16274 12114 16615 4 vdd
port 539 nsew
rlabel metal1 s 6606 15775 6642 16116 4 vdd
port 539 nsew
rlabel metal1 s 8334 14985 8370 15326 4 vdd
port 539 nsew
rlabel metal1 s 14574 11534 14610 11875 4 vdd
port 539 nsew
rlabel metal1 s 12078 23675 12114 24016 4 vdd
port 539 nsew
rlabel metal1 s 366 7875 402 8216 4 vdd
port 539 nsew
rlabel metal1 s 19086 21804 19122 22145 4 vdd
port 539 nsew
rlabel metal1 s 6606 8665 6642 9006 4 vdd
port 539 nsew
rlabel metal1 s 4110 14195 4146 14536 4 vdd
port 539 nsew
rlabel metal1 s 11598 17064 11634 17405 4 vdd
port 539 nsew
rlabel metal1 s 13326 1264 13362 1605 4 vdd
port 539 nsew
rlabel metal1 s 7854 22594 7890 22935 4 vdd
port 539 nsew
rlabel metal1 s 17838 24174 17874 24515 4 vdd
port 539 nsew
rlabel metal1 s 10830 24964 10866 25305 4 vdd
port 539 nsew
rlabel metal1 s 15342 5214 15378 5555 4 vdd
port 539 nsew
rlabel metal1 s 12078 3135 12114 3476 4 vdd
port 539 nsew
rlabel metal1 s 4590 14195 4626 14536 4 vdd
port 539 nsew
rlabel metal1 s 9102 474 9138 815 4 vdd
port 539 nsew
rlabel metal1 s 9102 12324 9138 12665 4 vdd
port 539 nsew
rlabel metal1 s 9102 7584 9138 7925 4 vdd
port 539 nsew
rlabel metal1 s 14094 24465 14130 24806 4 vdd
port 539 nsew
rlabel metal1 s 20334 24465 20370 24806 4 vdd
port 539 nsew
rlabel metal1 s 14574 23384 14610 23725 4 vdd
port 539 nsew
rlabel metal1 s 12078 21804 12114 22145 4 vdd
port 539 nsew
rlabel metal1 s 17070 1264 17106 1605 4 vdd
port 539 nsew
rlabel metal1 s 1614 21305 1650 21646 4 vdd
port 539 nsew
rlabel metal1 s 15822 6004 15858 6345 4 vdd
port 539 nsew
rlabel metal1 s 6606 7584 6642 7925 4 vdd
port 539 nsew
rlabel metal1 s 19086 6794 19122 7135 4 vdd
port 539 nsew
rlabel metal1 s 5838 14694 5874 15035 4 vdd
port 539 nsew
rlabel metal1 s 8334 1555 8370 1896 4 vdd
port 539 nsew
rlabel metal1 s 17838 19725 17874 20066 4 vdd
port 539 nsew
rlabel metal1 s 15822 18145 15858 18486 4 vdd
port 539 nsew
rlabel metal1 s 14094 10245 14130 10586 4 vdd
port 539 nsew
rlabel metal1 s 4110 21305 4146 21646 4 vdd
port 539 nsew
rlabel metal1 s 19566 17355 19602 17696 4 vdd
port 539 nsew
rlabel metal1 s 10350 17854 10386 18195 4 vdd
port 539 nsew
rlabel metal1 s 5838 19725 5874 20066 4 vdd
port 539 nsew
rlabel metal1 s 5358 23384 5394 23725 4 vdd
port 539 nsew
rlabel metal1 s 3342 9954 3378 10295 4 vdd
port 539 nsew
rlabel metal1 s 15822 22095 15858 22436 4 vdd
port 539 nsew
rlabel metal1 s 2094 14195 2130 14536 4 vdd
port 539 nsew
rlabel metal1 s 2094 18935 2130 19276 4 vdd
port 539 nsew
rlabel metal1 s 846 8374 882 8715 4 vdd
port 539 nsew
rlabel metal1 s 9582 22095 9618 22436 4 vdd
port 539 nsew
rlabel metal1 s 10830 25754 10866 26095 4 vdd
port 539 nsew
rlabel metal1 s 7854 21804 7890 22145 4 vdd
port 539 nsew
rlabel metal1 s 2094 20515 2130 20856 4 vdd
port 539 nsew
rlabel metal1 s 6606 1555 6642 1896 4 vdd
port 539 nsew
rlabel metal1 s 366 9455 402 9796 4 vdd
port 539 nsew
rlabel metal1 s 7854 1555 7890 1896 4 vdd
port 539 nsew
rlabel metal1 s 7854 17064 7890 17405 4 vdd
port 539 nsew
rlabel metal1 s 7086 2844 7122 3185 4 vdd
port 539 nsew
rlabel metal1 s 12078 474 12114 815 4 vdd
port 539 nsew
rlabel metal1 s 4110 11035 4146 11376 4 vdd
port 539 nsew
rlabel metal1 s 20334 14195 20370 14536 4 vdd
port 539 nsew
rlabel metal1 s 13326 18935 13362 19276 4 vdd
port 539 nsew
rlabel metal1 s 17070 15775 17106 16116 4 vdd
port 539 nsew
rlabel metal1 s 19566 18145 19602 18486 4 vdd
port 539 nsew
rlabel metal1 s 18318 2345 18354 2686 4 vdd
port 539 nsew
rlabel metal1 s 11598 20224 11634 20565 4 vdd
port 539 nsew
rlabel metal1 s 19086 14694 19122 15035 4 vdd
port 539 nsew
rlabel metal1 s 18318 9455 18354 9796 4 vdd
port 539 nsew
rlabel metal1 s 846 1555 882 1896 4 vdd
port 539 nsew
rlabel metal1 s 10350 1264 10386 1605 4 vdd
port 539 nsew
rlabel metal1 s 3342 24465 3378 24806 4 vdd
port 539 nsew
rlabel metal1 s 19566 7085 19602 7426 4 vdd
port 539 nsew
rlabel metal1 s 17070 25255 17106 25596 4 vdd
port 539 nsew
rlabel metal1 s 14574 474 14610 815 4 vdd
port 539 nsew
rlabel metal1 s 15342 23675 15378 24016 4 vdd
port 539 nsew
rlabel metal1 s 20334 17064 20370 17405 4 vdd
port 539 nsew
rlabel metal1 s 3342 24174 3378 24515 4 vdd
port 539 nsew
rlabel metal1 s 20334 7085 20370 7426 4 vdd
port 539 nsew
rlabel metal1 s 17838 11534 17874 11875 4 vdd
port 539 nsew
rlabel metal1 s 2094 765 2130 1106 4 vdd
port 539 nsew
rlabel metal1 s 7854 13904 7890 14245 4 vdd
port 539 nsew
rlabel metal1 s 19566 5505 19602 5846 4 vdd
port 539 nsew
rlabel metal1 s 13326 20515 13362 20856 4 vdd
port 539 nsew
rlabel metal1 s 4110 13904 4146 14245 4 vdd
port 539 nsew
rlabel metal1 s 10350 17355 10386 17696 4 vdd
port 539 nsew
rlabel metal1 s 2094 3925 2130 4266 4 vdd
port 539 nsew
rlabel metal1 s 4590 1555 4626 1896 4 vdd
port 539 nsew
rlabel metal1 s 19566 8374 19602 8715 4 vdd
port 539 nsew
rlabel metal1 s 18318 15775 18354 16116 4 vdd
port 539 nsew
rlabel metal1 s 2862 21804 2898 22145 4 vdd
port 539 nsew
rlabel metal1 s 10830 9455 10866 9796 4 vdd
port 539 nsew
rlabel metal1 s 10350 22095 10386 22436 4 vdd
port 539 nsew
rlabel metal1 s 20334 12615 20370 12956 4 vdd
port 539 nsew
rlabel metal1 s 14094 18644 14130 18985 4 vdd
port 539 nsew
rlabel metal1 s 12846 9455 12882 9796 4 vdd
port 539 nsew
rlabel metal1 s 15342 13405 15378 13746 4 vdd
port 539 nsew
rlabel metal1 s 9582 10245 9618 10586 4 vdd
port 539 nsew
rlabel metal1 s 3342 16274 3378 16615 4 vdd
port 539 nsew
rlabel metal1 s 366 11825 402 12166 4 vdd
port 539 nsew
rlabel metal1 s 20334 14985 20370 15326 4 vdd
port 539 nsew
rlabel metal1 s 20814 20224 20850 20565 4 vdd
port 539 nsew
rlabel metal1 s 7086 1555 7122 1896 4 vdd
port 539 nsew
rlabel metal1 s 2094 7584 2130 7925 4 vdd
port 539 nsew
rlabel metal1 s 19086 21014 19122 21355 4 vdd
port 539 nsew
rlabel metal1 s 15822 22594 15858 22935 4 vdd
port 539 nsew
rlabel metal1 s 14094 24174 14130 24515 4 vdd
port 539 nsew
rlabel metal1 s 2094 9455 2130 9796 4 vdd
port 539 nsew
rlabel metal1 s 9582 6004 9618 6345 4 vdd
port 539 nsew
rlabel metal1 s 17070 8374 17106 8715 4 vdd
port 539 nsew
rlabel metal1 s 10830 16565 10866 16906 4 vdd
port 539 nsew
rlabel metal1 s 16590 20515 16626 20856 4 vdd
port 539 nsew
rlabel metal1 s 2862 23675 2898 24016 4 vdd
port 539 nsew
rlabel metal1 s 17838 16274 17874 16615 4 vdd
port 539 nsew
rlabel metal1 s 19086 15484 19122 15825 4 vdd
port 539 nsew
rlabel metal1 s 366 8374 402 8715 4 vdd
port 539 nsew
rlabel metal1 s 5358 14985 5394 15326 4 vdd
port 539 nsew
rlabel metal1 s 12078 11534 12114 11875 4 vdd
port 539 nsew
rlabel metal1 s 1614 10245 1650 10586 4 vdd
port 539 nsew
rlabel metal1 s 8334 22885 8370 23226 4 vdd
port 539 nsew
rlabel metal1 s 12078 24465 12114 24806 4 vdd
port 539 nsew
rlabel metal1 s 1614 5505 1650 5846 4 vdd
port 539 nsew
rlabel metal1 s 17070 4424 17106 4765 4 vdd
port 539 nsew
rlabel metal1 s 3342 765 3378 1106 4 vdd
port 539 nsew
rlabel metal1 s 9102 23384 9138 23725 4 vdd
port 539 nsew
rlabel metal1 s 2862 12615 2898 12956 4 vdd
port 539 nsew
rlabel metal1 s 19086 24465 19122 24806 4 vdd
port 539 nsew
rlabel metal1 s 1614 8665 1650 9006 4 vdd
port 539 nsew
rlabel metal1 s 19566 765 19602 1106 4 vdd
port 539 nsew
rlabel metal1 s 17070 13904 17106 14245 4 vdd
port 539 nsew
rlabel metal1 s 13326 14694 13362 15035 4 vdd
port 539 nsew
rlabel metal1 s 9102 24465 9138 24806 4 vdd
port 539 nsew
rlabel metal1 s 17838 2844 17874 3185 4 vdd
port 539 nsew
rlabel metal1 s 18318 24964 18354 25305 4 vdd
port 539 nsew
rlabel metal1 s 9582 23675 9618 24016 4 vdd
port 539 nsew
rlabel metal1 s 2094 16274 2130 16615 4 vdd
port 539 nsew
rlabel metal1 s 14574 10245 14610 10586 4 vdd
port 539 nsew
rlabel metal1 s 15342 18935 15378 19276 4 vdd
port 539 nsew
rlabel metal1 s 13326 18644 13362 18985 4 vdd
port 539 nsew
rlabel metal1 s 14094 8665 14130 9006 4 vdd
port 539 nsew
rlabel metal1 s 8334 6004 8370 6345 4 vdd
port 539 nsew
rlabel metal1 s 19086 4424 19122 4765 4 vdd
port 539 nsew
rlabel metal1 s 5358 15484 5394 15825 4 vdd
port 539 nsew
rlabel metal1 s 3342 15484 3378 15825 4 vdd
port 539 nsew
rlabel metal1 s 366 15775 402 16116 4 vdd
port 539 nsew
rlabel metal1 s 8334 24465 8370 24806 4 vdd
port 539 nsew
rlabel metal1 s 846 9954 882 10295 4 vdd
port 539 nsew
rlabel metal1 s 4590 3135 4626 3476 4 vdd
port 539 nsew
rlabel metal1 s 13326 23675 13362 24016 4 vdd
port 539 nsew
rlabel metal1 s 9102 9164 9138 9505 4 vdd
port 539 nsew
rlabel metal1 s 846 -25 882 316 4 vdd
port 539 nsew
rlabel metal1 s 7086 1264 7122 1605 4 vdd
port 539 nsew
rlabel metal1 s 2862 14985 2898 15326 4 vdd
port 539 nsew
rlabel metal1 s 11598 23675 11634 24016 4 vdd
port 539 nsew
rlabel metal1 s 4110 6794 4146 7135 4 vdd
port 539 nsew
rlabel metal1 s 11598 11035 11634 11376 4 vdd
port 539 nsew
rlabel metal1 s 6606 3634 6642 3975 4 vdd
port 539 nsew
rlabel metal1 s 6606 13405 6642 13746 4 vdd
port 539 nsew
rlabel metal1 s 9582 12324 9618 12665 4 vdd
port 539 nsew
rlabel metal1 s 9102 23675 9138 24016 4 vdd
port 539 nsew
rlabel metal1 s 20814 18145 20850 18486 4 vdd
port 539 nsew
rlabel metal1 s 9102 15775 9138 16116 4 vdd
port 539 nsew
rlabel metal1 s 17070 4715 17106 5056 4 vdd
port 539 nsew
rlabel metal1 s 4590 474 4626 815 4 vdd
port 539 nsew
rlabel metal1 s 3342 20224 3378 20565 4 vdd
port 539 nsew
rlabel metal1 s 13326 24964 13362 25305 4 vdd
port 539 nsew
rlabel metal1 s 17838 21305 17874 21646 4 vdd
port 539 nsew
rlabel metal1 s 20334 -25 20370 316 4 vdd
port 539 nsew
rlabel metal1 s 17838 20224 17874 20565 4 vdd
port 539 nsew
rlabel metal1 s 12846 3925 12882 4266 4 vdd
port 539 nsew
rlabel metal1 s 5358 19434 5394 19775 4 vdd
port 539 nsew
rlabel metal1 s 18318 18145 18354 18486 4 vdd
port 539 nsew
rlabel metal1 s 9582 9164 9618 9505 4 vdd
port 539 nsew
rlabel metal1 s 11598 19725 11634 20066 4 vdd
port 539 nsew
rlabel metal1 s 5838 20515 5874 20856 4 vdd
port 539 nsew
rlabel metal1 s 3342 25255 3378 25596 4 vdd
port 539 nsew
rlabel metal1 s 11598 1555 11634 1896 4 vdd
port 539 nsew
rlabel metal1 s 14574 22885 14610 23226 4 vdd
port 539 nsew
rlabel metal1 s 12078 15484 12114 15825 4 vdd
port 539 nsew
rlabel metal1 s 1614 24465 1650 24806 4 vdd
port 539 nsew
rlabel metal1 s 19566 6004 19602 6345 4 vdd
port 539 nsew
rlabel metal1 s 6606 -25 6642 316 4 vdd
port 539 nsew
rlabel metal1 s 17070 11534 17106 11875 4 vdd
port 539 nsew
rlabel metal1 s 14094 9164 14130 9505 4 vdd
port 539 nsew
rlabel metal1 s 11598 14985 11634 15326 4 vdd
port 539 nsew
rlabel metal1 s 12846 21014 12882 21355 4 vdd
port 539 nsew
rlabel metal1 s 19086 5214 19122 5555 4 vdd
port 539 nsew
rlabel metal1 s 18318 11035 18354 11376 4 vdd
port 539 nsew
rlabel metal1 s 4590 20224 4626 20565 4 vdd
port 539 nsew
rlabel metal1 s 14094 11534 14130 11875 4 vdd
port 539 nsew
rlabel metal1 s 17838 3925 17874 4266 4 vdd
port 539 nsew
rlabel metal1 s 20814 7875 20850 8216 4 vdd
port 539 nsew
rlabel metal1 s 18318 2054 18354 2395 4 vdd
port 539 nsew
rlabel metal1 s 20334 4715 20370 5056 4 vdd
port 539 nsew
rlabel metal1 s 12078 8665 12114 9006 4 vdd
port 539 nsew
rlabel metal1 s 15822 11035 15858 11376 4 vdd
port 539 nsew
rlabel metal1 s 10830 6295 10866 6636 4 vdd
port 539 nsew
rlabel metal1 s 12078 6004 12114 6345 4 vdd
port 539 nsew
rlabel metal1 s 10350 15484 10386 15825 4 vdd
port 539 nsew
rlabel metal1 s 12078 14694 12114 15035 4 vdd
port 539 nsew
rlabel metal1 s 15822 17854 15858 18195 4 vdd
port 539 nsew
rlabel metal1 s 7086 5505 7122 5846 4 vdd
port 539 nsew
rlabel metal1 s 366 18644 402 18985 4 vdd
port 539 nsew
rlabel metal1 s 10350 8374 10386 8715 4 vdd
port 539 nsew
rlabel metal1 s 18318 5505 18354 5846 4 vdd
port 539 nsew
rlabel metal1 s 17838 22885 17874 23226 4 vdd
port 539 nsew
rlabel metal1 s 19566 24174 19602 24515 4 vdd
port 539 nsew
rlabel metal1 s 19566 15484 19602 15825 4 vdd
port 539 nsew
rlabel metal1 s 15342 22095 15378 22436 4 vdd
port 539 nsew
rlabel metal1 s 1614 9455 1650 9796 4 vdd
port 539 nsew
rlabel metal1 s 9582 18644 9618 18985 4 vdd
port 539 nsew
rlabel metal1 s 7086 9954 7122 10295 4 vdd
port 539 nsew
rlabel metal1 s 13326 -25 13362 316 4 vdd
port 539 nsew
rlabel metal1 s 3342 -25 3378 316 4 vdd
port 539 nsew
rlabel metal1 s 846 15484 882 15825 4 vdd
port 539 nsew
rlabel metal1 s 17838 765 17874 1106 4 vdd
port 539 nsew
rlabel metal1 s 4110 6295 4146 6636 4 vdd
port 539 nsew
rlabel metal1 s 5358 -25 5394 316 4 vdd
port 539 nsew
rlabel metal1 s 10350 11035 10386 11376 4 vdd
port 539 nsew
rlabel metal1 s 7086 21305 7122 21646 4 vdd
port 539 nsew
rlabel metal1 s 12078 12615 12114 12956 4 vdd
port 539 nsew
rlabel metal1 s 9582 13904 9618 14245 4 vdd
port 539 nsew
rlabel metal1 s 2862 17064 2898 17405 4 vdd
port 539 nsew
rlabel metal1 s 18318 21804 18354 22145 4 vdd
port 539 nsew
rlabel metal1 s 20814 14985 20850 15326 4 vdd
port 539 nsew
rlabel metal1 s 17838 14195 17874 14536 4 vdd
port 539 nsew
rlabel metal1 s 6606 22095 6642 22436 4 vdd
port 539 nsew
rlabel metal1 s 12846 24465 12882 24806 4 vdd
port 539 nsew
rlabel metal1 s 366 6794 402 7135 4 vdd
port 539 nsew
rlabel metal1 s 16590 21014 16626 21355 4 vdd
port 539 nsew
rlabel metal1 s 9102 20224 9138 20565 4 vdd
port 539 nsew
rlabel metal1 s 2094 20224 2130 20565 4 vdd
port 539 nsew
rlabel metal1 s 19566 25754 19602 26095 4 vdd
port 539 nsew
rlabel metal1 s 19566 8665 19602 9006 4 vdd
port 539 nsew
rlabel metal1 s 7086 15775 7122 16116 4 vdd
port 539 nsew
rlabel metal1 s 4110 765 4146 1106 4 vdd
port 539 nsew
rlabel metal1 s 5838 13405 5874 13746 4 vdd
port 539 nsew
rlabel metal1 s 5838 2054 5874 2395 4 vdd
port 539 nsew
rlabel metal1 s 7854 18935 7890 19276 4 vdd
port 539 nsew
rlabel metal1 s 3342 9455 3378 9796 4 vdd
port 539 nsew
rlabel metal1 s 18318 474 18354 815 4 vdd
port 539 nsew
rlabel metal1 s 14574 13904 14610 14245 4 vdd
port 539 nsew
rlabel metal1 s 366 11035 402 11376 4 vdd
port 539 nsew
rlabel metal1 s 10350 18935 10386 19276 4 vdd
port 539 nsew
rlabel metal1 s 4110 11534 4146 11875 4 vdd
port 539 nsew
rlabel metal1 s 10350 765 10386 1106 4 vdd
port 539 nsew
rlabel metal1 s 19086 8374 19122 8715 4 vdd
port 539 nsew
rlabel metal1 s 15822 24964 15858 25305 4 vdd
port 539 nsew
rlabel metal1 s 13326 22095 13362 22436 4 vdd
port 539 nsew
rlabel metal1 s 18318 24174 18354 24515 4 vdd
port 539 nsew
rlabel metal1 s 7086 22594 7122 22935 4 vdd
port 539 nsew
rlabel metal1 s 2862 9954 2898 10295 4 vdd
port 539 nsew
rlabel metal1 s 20814 3135 20850 3476 4 vdd
port 539 nsew
rlabel metal1 s 1614 4424 1650 4765 4 vdd
port 539 nsew
rlabel metal1 s 18318 14694 18354 15035 4 vdd
port 539 nsew
rlabel metal1 s 15822 14195 15858 14536 4 vdd
port 539 nsew
rlabel metal1 s 11598 7085 11634 7426 4 vdd
port 539 nsew
rlabel metal1 s 3342 15775 3378 16116 4 vdd
port 539 nsew
rlabel metal1 s 5358 24964 5394 25305 4 vdd
port 539 nsew
rlabel metal1 s 7854 9455 7890 9796 4 vdd
port 539 nsew
rlabel metal1 s 6606 15484 6642 15825 4 vdd
port 539 nsew
rlabel metal1 s 5358 8374 5394 8715 4 vdd
port 539 nsew
rlabel metal1 s 15822 5505 15858 5846 4 vdd
port 539 nsew
rlabel metal1 s 4590 21014 4626 21355 4 vdd
port 539 nsew
rlabel metal1 s 20814 3634 20850 3975 4 vdd
port 539 nsew
rlabel metal1 s 7854 14985 7890 15326 4 vdd
port 539 nsew
rlabel metal1 s 846 5214 882 5555 4 vdd
port 539 nsew
rlabel metal1 s 17838 3135 17874 3476 4 vdd
port 539 nsew
rlabel metal1 s 20334 18935 20370 19276 4 vdd
port 539 nsew
rlabel metal1 s 2862 25255 2898 25596 4 vdd
port 539 nsew
rlabel metal1 s 10830 7584 10866 7925 4 vdd
port 539 nsew
rlabel metal1 s 20334 18145 20370 18486 4 vdd
port 539 nsew
rlabel metal1 s 4590 17854 4626 18195 4 vdd
port 539 nsew
rlabel metal1 s 15822 11534 15858 11875 4 vdd
port 539 nsew
rlabel metal1 s 10350 21804 10386 22145 4 vdd
port 539 nsew
rlabel metal1 s 7854 474 7890 815 4 vdd
port 539 nsew
rlabel metal1 s 12846 14985 12882 15326 4 vdd
port 539 nsew
rlabel metal1 s 14574 6004 14610 6345 4 vdd
port 539 nsew
rlabel metal1 s 5838 15775 5874 16116 4 vdd
port 539 nsew
rlabel metal1 s 3342 22594 3378 22935 4 vdd
port 539 nsew
rlabel metal1 s 5838 3925 5874 4266 4 vdd
port 539 nsew
rlabel metal1 s 4590 2054 4626 2395 4 vdd
port 539 nsew
rlabel metal1 s 12846 5505 12882 5846 4 vdd
port 539 nsew
rlabel metal1 s 18318 4424 18354 4765 4 vdd
port 539 nsew
rlabel metal1 s 9582 2345 9618 2686 4 vdd
port 539 nsew
rlabel metal1 s 6606 16565 6642 16906 4 vdd
port 539 nsew
rlabel metal1 s 10350 22885 10386 23226 4 vdd
port 539 nsew
rlabel metal1 s 2862 8665 2898 9006 4 vdd
port 539 nsew
rlabel metal1 s 4590 21804 4626 22145 4 vdd
port 539 nsew
rlabel metal1 s 7854 22095 7890 22436 4 vdd
port 539 nsew
rlabel metal1 s 20334 14694 20370 15035 4 vdd
port 539 nsew
rlabel metal1 s 17838 1555 17874 1896 4 vdd
port 539 nsew
rlabel metal1 s 15822 13114 15858 13455 4 vdd
port 539 nsew
rlabel metal1 s 4590 10245 4626 10586 4 vdd
port 539 nsew
rlabel metal1 s 10830 5214 10866 5555 4 vdd
port 539 nsew
rlabel metal1 s 10350 4715 10386 5056 4 vdd
port 539 nsew
rlabel metal1 s 4110 25255 4146 25596 4 vdd
port 539 nsew
rlabel metal1 s 846 22594 882 22935 4 vdd
port 539 nsew
rlabel metal1 s 2862 16565 2898 16906 4 vdd
port 539 nsew
rlabel metal1 s 2094 14694 2130 15035 4 vdd
port 539 nsew
rlabel metal1 s 8334 18644 8370 18985 4 vdd
port 539 nsew
rlabel metal1 s 846 14694 882 15035 4 vdd
port 539 nsew
rlabel metal1 s 14094 12615 14130 12956 4 vdd
port 539 nsew
rlabel metal1 s 4110 12324 4146 12665 4 vdd
port 539 nsew
rlabel metal1 s 20334 4424 20370 4765 4 vdd
port 539 nsew
rlabel metal1 s 13326 9954 13362 10295 4 vdd
port 539 nsew
rlabel metal1 s 17070 19725 17106 20066 4 vdd
port 539 nsew
rlabel metal1 s 846 19434 882 19775 4 vdd
port 539 nsew
rlabel metal1 s 12846 24174 12882 24515 4 vdd
port 539 nsew
rlabel metal1 s 14574 7875 14610 8216 4 vdd
port 539 nsew
rlabel metal1 s 4590 25754 4626 26095 4 vdd
port 539 nsew
rlabel metal1 s 14094 19725 14130 20066 4 vdd
port 539 nsew
rlabel metal1 s 9582 21014 9618 21355 4 vdd
port 539 nsew
rlabel metal1 s 11598 6295 11634 6636 4 vdd
port 539 nsew
rlabel metal1 s 1614 3634 1650 3975 4 vdd
port 539 nsew
rlabel metal1 s 10350 13114 10386 13455 4 vdd
port 539 nsew
rlabel metal1 s 5838 2844 5874 3185 4 vdd
port 539 nsew
rlabel metal1 s 10830 17355 10866 17696 4 vdd
port 539 nsew
rlabel metal1 s 1614 2345 1650 2686 4 vdd
port 539 nsew
rlabel metal1 s 18318 20224 18354 20565 4 vdd
port 539 nsew
rlabel metal1 s 4110 2345 4146 2686 4 vdd
port 539 nsew
rlabel metal1 s 13326 21014 13362 21355 4 vdd
port 539 nsew
rlabel metal1 s 2094 25754 2130 26095 4 vdd
port 539 nsew
rlabel metal1 s 7854 -25 7890 316 4 vdd
port 539 nsew
rlabel metal1 s 14574 23675 14610 24016 4 vdd
port 539 nsew
rlabel metal1 s 7854 4715 7890 5056 4 vdd
port 539 nsew
rlabel metal1 s 17070 9164 17106 9505 4 vdd
port 539 nsew
rlabel metal1 s 4110 474 4146 815 4 vdd
port 539 nsew
rlabel metal1 s 9582 14985 9618 15326 4 vdd
port 539 nsew
rlabel metal1 s 11598 21014 11634 21355 4 vdd
port 539 nsew
rlabel metal1 s 6606 6004 6642 6345 4 vdd
port 539 nsew
rlabel metal1 s 8334 -25 8370 316 4 vdd
port 539 nsew
rlabel metal1 s 19566 19434 19602 19775 4 vdd
port 539 nsew
rlabel metal1 s 12078 13114 12114 13455 4 vdd
port 539 nsew
rlabel metal1 s 366 24964 402 25305 4 vdd
port 539 nsew
rlabel metal1 s 3342 14985 3378 15326 4 vdd
port 539 nsew
rlabel metal1 s 15342 15484 15378 15825 4 vdd
port 539 nsew
rlabel metal1 s 14094 8374 14130 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 10744 9138 11085 4 vdd
port 539 nsew
rlabel metal1 s 16590 17064 16626 17405 4 vdd
port 539 nsew
rlabel metal1 s 19086 2345 19122 2686 4 vdd
port 539 nsew
rlabel metal1 s 19566 12324 19602 12665 4 vdd
port 539 nsew
rlabel metal1 s 6606 5505 6642 5846 4 vdd
port 539 nsew
rlabel metal1 s 7854 3634 7890 3975 4 vdd
port 539 nsew
rlabel metal1 s 4110 10245 4146 10586 4 vdd
port 539 nsew
rlabel metal1 s 20334 23384 20370 23725 4 vdd
port 539 nsew
rlabel metal1 s 3342 3135 3378 3476 4 vdd
port 539 nsew
rlabel metal1 s 7086 6004 7122 6345 4 vdd
port 539 nsew
rlabel metal1 s 14574 19725 14610 20066 4 vdd
port 539 nsew
rlabel metal1 s 7086 3925 7122 4266 4 vdd
port 539 nsew
rlabel metal1 s 20334 765 20370 1106 4 vdd
port 539 nsew
rlabel metal1 s 19566 14195 19602 14536 4 vdd
port 539 nsew
rlabel metal1 s 9102 22594 9138 22935 4 vdd
port 539 nsew
rlabel metal1 s 20814 5214 20850 5555 4 vdd
port 539 nsew
rlabel metal1 s 12846 20515 12882 20856 4 vdd
port 539 nsew
rlabel metal1 s 1614 18644 1650 18985 4 vdd
port 539 nsew
rlabel metal1 s 2094 7085 2130 7426 4 vdd
port 539 nsew
rlabel metal1 s 5358 14694 5394 15035 4 vdd
port 539 nsew
rlabel metal1 s 15342 765 15378 1106 4 vdd
port 539 nsew
rlabel metal1 s 14094 3135 14130 3476 4 vdd
port 539 nsew
rlabel metal1 s 9582 7085 9618 7426 4 vdd
port 539 nsew
rlabel metal1 s 20334 2345 20370 2686 4 vdd
port 539 nsew
rlabel metal1 s 10830 6794 10866 7135 4 vdd
port 539 nsew
rlabel metal1 s 19566 22885 19602 23226 4 vdd
port 539 nsew
rlabel metal1 s 14094 17064 14130 17405 4 vdd
port 539 nsew
rlabel metal1 s 16590 15484 16626 15825 4 vdd
port 539 nsew
rlabel metal1 s 4110 17854 4146 18195 4 vdd
port 539 nsew
rlabel metal1 s 13326 19725 13362 20066 4 vdd
port 539 nsew
rlabel metal1 s 6606 21014 6642 21355 4 vdd
port 539 nsew
rlabel metal1 s 17070 9954 17106 10295 4 vdd
port 539 nsew
rlabel metal1 s 15822 7085 15858 7426 4 vdd
port 539 nsew
rlabel metal1 s 3342 17064 3378 17405 4 vdd
port 539 nsew
rlabel metal1 s 8334 7875 8370 8216 4 vdd
port 539 nsew
rlabel metal1 s 1614 14195 1650 14536 4 vdd
port 539 nsew
rlabel metal1 s 366 5505 402 5846 4 vdd
port 539 nsew
rlabel metal1 s 4110 21014 4146 21355 4 vdd
port 539 nsew
rlabel metal1 s 15822 25754 15858 26095 4 vdd
port 539 nsew
rlabel metal1 s 5358 10744 5394 11085 4 vdd
port 539 nsew
rlabel metal1 s 5358 474 5394 815 4 vdd
port 539 nsew
rlabel metal1 s 6606 20515 6642 20856 4 vdd
port 539 nsew
rlabel metal1 s 366 23384 402 23725 4 vdd
port 539 nsew
rlabel metal1 s 5358 8665 5394 9006 4 vdd
port 539 nsew
rlabel metal1 s 9102 6295 9138 6636 4 vdd
port 539 nsew
rlabel metal1 s 4110 22885 4146 23226 4 vdd
port 539 nsew
rlabel metal1 s 19086 16565 19122 16906 4 vdd
port 539 nsew
rlabel metal1 s 13326 17355 13362 17696 4 vdd
port 539 nsew
rlabel metal1 s 6606 23675 6642 24016 4 vdd
port 539 nsew
rlabel metal1 s 846 19725 882 20066 4 vdd
port 539 nsew
rlabel metal1 s 4590 5505 4626 5846 4 vdd
port 539 nsew
rlabel metal1 s 9102 25255 9138 25596 4 vdd
port 539 nsew
rlabel metal1 s 15342 2054 15378 2395 4 vdd
port 539 nsew
rlabel metal1 s 10350 19725 10386 20066 4 vdd
port 539 nsew
rlabel metal1 s 19566 3634 19602 3975 4 vdd
port 539 nsew
rlabel metal1 s 13326 3634 13362 3975 4 vdd
port 539 nsew
rlabel metal1 s 10350 25255 10386 25596 4 vdd
port 539 nsew
rlabel metal1 s 18318 9164 18354 9505 4 vdd
port 539 nsew
rlabel metal1 s 7854 6004 7890 6345 4 vdd
port 539 nsew
rlabel metal1 s 3342 11825 3378 12166 4 vdd
port 539 nsew
rlabel metal1 s 11598 15775 11634 16116 4 vdd
port 539 nsew
rlabel metal1 s 20334 19725 20370 20066 4 vdd
port 539 nsew
rlabel metal1 s 12078 22885 12114 23226 4 vdd
port 539 nsew
rlabel metal1 s 10830 22594 10866 22935 4 vdd
port 539 nsew
rlabel metal1 s 10350 25754 10386 26095 4 vdd
port 539 nsew
rlabel metal1 s 14574 25754 14610 26095 4 vdd
port 539 nsew
rlabel metal1 s 19566 23384 19602 23725 4 vdd
port 539 nsew
rlabel metal1 s 5358 21014 5394 21355 4 vdd
port 539 nsew
rlabel metal1 s 10350 20515 10386 20856 4 vdd
port 539 nsew
rlabel metal1 s 2094 8665 2130 9006 4 vdd
port 539 nsew
rlabel metal1 s 12078 1264 12114 1605 4 vdd
port 539 nsew
rlabel metal1 s 15342 6794 15378 7135 4 vdd
port 539 nsew
rlabel metal1 s 19086 13904 19122 14245 4 vdd
port 539 nsew
rlabel metal1 s 11598 1264 11634 1605 4 vdd
port 539 nsew
rlabel metal1 s 11598 17355 11634 17696 4 vdd
port 539 nsew
rlabel metal1 s 9582 24964 9618 25305 4 vdd
port 539 nsew
rlabel metal1 s 16590 21804 16626 22145 4 vdd
port 539 nsew
rlabel metal1 s 7086 765 7122 1106 4 vdd
port 539 nsew
rlabel metal1 s 10350 11825 10386 12166 4 vdd
port 539 nsew
rlabel metal1 s 12846 13114 12882 13455 4 vdd
port 539 nsew
rlabel metal1 s 20814 20515 20850 20856 4 vdd
port 539 nsew
rlabel metal1 s 17838 8374 17874 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 17854 9138 18195 4 vdd
port 539 nsew
rlabel metal1 s 9582 21804 9618 22145 4 vdd
port 539 nsew
rlabel metal1 s 10830 11534 10866 11875 4 vdd
port 539 nsew
rlabel metal1 s 17070 13114 17106 13455 4 vdd
port 539 nsew
rlabel metal1 s 14094 12324 14130 12665 4 vdd
port 539 nsew
rlabel metal1 s 8334 15775 8370 16116 4 vdd
port 539 nsew
rlabel metal1 s 366 4715 402 5056 4 vdd
port 539 nsew
rlabel metal1 s 20814 14195 20850 14536 4 vdd
port 539 nsew
rlabel metal1 s 12078 14195 12114 14536 4 vdd
port 539 nsew
rlabel metal1 s 9102 3925 9138 4266 4 vdd
port 539 nsew
rlabel metal1 s 2862 4424 2898 4765 4 vdd
port 539 nsew
rlabel metal1 s 20334 5214 20370 5555 4 vdd
port 539 nsew
rlabel metal1 s 7854 19434 7890 19775 4 vdd
port 539 nsew
rlabel metal1 s 19566 23675 19602 24016 4 vdd
port 539 nsew
rlabel metal1 s 846 2844 882 3185 4 vdd
port 539 nsew
rlabel metal1 s 2094 24964 2130 25305 4 vdd
port 539 nsew
rlabel metal1 s 4110 4424 4146 4765 4 vdd
port 539 nsew
rlabel metal1 s 9102 8665 9138 9006 4 vdd
port 539 nsew
rlabel metal1 s 9102 5214 9138 5555 4 vdd
port 539 nsew
rlabel metal1 s 19566 11825 19602 12166 4 vdd
port 539 nsew
rlabel metal1 s 366 10744 402 11085 4 vdd
port 539 nsew
rlabel metal1 s 2094 18644 2130 18985 4 vdd
port 539 nsew
rlabel metal1 s 7086 6794 7122 7135 4 vdd
port 539 nsew
rlabel metal1 s 17838 9455 17874 9796 4 vdd
port 539 nsew
rlabel metal1 s 10830 3634 10866 3975 4 vdd
port 539 nsew
rlabel metal1 s 10830 17064 10866 17405 4 vdd
port 539 nsew
rlabel metal1 s 10350 12324 10386 12665 4 vdd
port 539 nsew
rlabel metal1 s 17070 22095 17106 22436 4 vdd
port 539 nsew
rlabel metal1 s 16590 25255 16626 25596 4 vdd
port 539 nsew
rlabel metal1 s 5838 1264 5874 1605 4 vdd
port 539 nsew
rlabel metal1 s 14094 2054 14130 2395 4 vdd
port 539 nsew
rlabel metal1 s 6606 13904 6642 14245 4 vdd
port 539 nsew
rlabel metal1 s 16590 19725 16626 20066 4 vdd
port 539 nsew
rlabel metal1 s 10830 1555 10866 1896 4 vdd
port 539 nsew
rlabel metal1 s 3342 11534 3378 11875 4 vdd
port 539 nsew
rlabel metal1 s 3342 24964 3378 25305 4 vdd
port 539 nsew
rlabel metal1 s 16590 765 16626 1106 4 vdd
port 539 nsew
rlabel metal1 s 17838 2054 17874 2395 4 vdd
port 539 nsew
rlabel metal1 s 12078 10245 12114 10586 4 vdd
port 539 nsew
rlabel metal1 s 10350 13405 10386 13746 4 vdd
port 539 nsew
rlabel metal1 s 12846 4715 12882 5056 4 vdd
port 539 nsew
rlabel metal1 s 12846 15775 12882 16116 4 vdd
port 539 nsew
rlabel metal1 s 8334 6794 8370 7135 4 vdd
port 539 nsew
rlabel metal1 s 2862 7584 2898 7925 4 vdd
port 539 nsew
rlabel metal1 s 17838 8665 17874 9006 4 vdd
port 539 nsew
rlabel metal1 s 2862 5214 2898 5555 4 vdd
port 539 nsew
rlabel metal1 s 10830 9954 10866 10295 4 vdd
port 539 nsew
rlabel metal1 s 18318 14985 18354 15326 4 vdd
port 539 nsew
rlabel metal1 s 5358 4424 5394 4765 4 vdd
port 539 nsew
rlabel metal1 s 5838 -25 5874 316 4 vdd
port 539 nsew
rlabel metal1 s 12078 18644 12114 18985 4 vdd
port 539 nsew
rlabel metal1 s 1614 7875 1650 8216 4 vdd
port 539 nsew
rlabel metal1 s 20814 10245 20850 10586 4 vdd
port 539 nsew
rlabel metal1 s 7086 11035 7122 11376 4 vdd
port 539 nsew
rlabel metal1 s 14574 9954 14610 10295 4 vdd
port 539 nsew
rlabel metal1 s 16590 14195 16626 14536 4 vdd
port 539 nsew
rlabel metal1 s 1614 14985 1650 15326 4 vdd
port 539 nsew
rlabel metal1 s 13326 19434 13362 19775 4 vdd
port 539 nsew
rlabel metal1 s 10830 20224 10866 20565 4 vdd
port 539 nsew
rlabel metal1 s 7086 18935 7122 19276 4 vdd
port 539 nsew
rlabel metal1 s 12846 8374 12882 8715 4 vdd
port 539 nsew
rlabel metal1 s 9102 10245 9138 10586 4 vdd
port 539 nsew
rlabel metal1 s 5838 6004 5874 6345 4 vdd
port 539 nsew
rlabel metal1 s 17838 22095 17874 22436 4 vdd
port 539 nsew
rlabel metal1 s 4590 24174 4626 24515 4 vdd
port 539 nsew
rlabel metal1 s 15822 24465 15858 24806 4 vdd
port 539 nsew
rlabel metal1 s 12846 23384 12882 23725 4 vdd
port 539 nsew
rlabel metal1 s 10350 474 10386 815 4 vdd
port 539 nsew
rlabel metal1 s 14094 7584 14130 7925 4 vdd
port 539 nsew
rlabel metal1 s 10830 7875 10866 8216 4 vdd
port 539 nsew
rlabel metal1 s 10830 18145 10866 18486 4 vdd
port 539 nsew
rlabel metal1 s 10830 20515 10866 20856 4 vdd
port 539 nsew
rlabel metal1 s 10830 3925 10866 4266 4 vdd
port 539 nsew
rlabel metal1 s 20814 474 20850 815 4 vdd
port 539 nsew
rlabel metal1 s 14574 22095 14610 22436 4 vdd
port 539 nsew
rlabel metal1 s 20334 16274 20370 16615 4 vdd
port 539 nsew
rlabel metal1 s 12846 17064 12882 17405 4 vdd
port 539 nsew
rlabel metal1 s 20334 15775 20370 16116 4 vdd
port 539 nsew
rlabel metal1 s 5838 24964 5874 25305 4 vdd
port 539 nsew
rlabel metal1 s 10830 14694 10866 15035 4 vdd
port 539 nsew
rlabel metal1 s 3342 2844 3378 3185 4 vdd
port 539 nsew
rlabel metal1 s 13326 14195 13362 14536 4 vdd
port 539 nsew
rlabel metal1 s 846 6295 882 6636 4 vdd
port 539 nsew
rlabel metal1 s 846 6004 882 6345 4 vdd
port 539 nsew
rlabel metal1 s 8334 23675 8370 24016 4 vdd
port 539 nsew
rlabel metal1 s 14574 13405 14610 13746 4 vdd
port 539 nsew
rlabel metal1 s 18318 12615 18354 12956 4 vdd
port 539 nsew
rlabel metal1 s 6606 20224 6642 20565 4 vdd
port 539 nsew
rlabel metal1 s 19566 9164 19602 9505 4 vdd
port 539 nsew
rlabel metal1 s 20334 11825 20370 12166 4 vdd
port 539 nsew
rlabel metal1 s 14094 13405 14130 13746 4 vdd
port 539 nsew
rlabel metal1 s 4590 6004 4626 6345 4 vdd
port 539 nsew
rlabel metal1 s 846 15775 882 16116 4 vdd
port 539 nsew
rlabel metal1 s 10830 17854 10866 18195 4 vdd
port 539 nsew
rlabel metal1 s 10830 19434 10866 19775 4 vdd
port 539 nsew
rlabel metal1 s 17070 2345 17106 2686 4 vdd
port 539 nsew
rlabel metal1 s 17070 18644 17106 18985 4 vdd
port 539 nsew
rlabel metal1 s 16590 5505 16626 5846 4 vdd
port 539 nsew
rlabel metal1 s 7086 20224 7122 20565 4 vdd
port 539 nsew
rlabel metal1 s 5838 14195 5874 14536 4 vdd
port 539 nsew
rlabel metal1 s 15342 22594 15378 22935 4 vdd
port 539 nsew
rlabel metal1 s 17838 15775 17874 16116 4 vdd
port 539 nsew
rlabel metal1 s 10830 14195 10866 14536 4 vdd
port 539 nsew
rlabel metal1 s 20334 7584 20370 7925 4 vdd
port 539 nsew
rlabel metal1 s 14574 2844 14610 3185 4 vdd
port 539 nsew
rlabel metal1 s 13326 11825 13362 12166 4 vdd
port 539 nsew
rlabel metal1 s 17838 4424 17874 4765 4 vdd
port 539 nsew
rlabel metal1 s 8334 23384 8370 23725 4 vdd
port 539 nsew
rlabel metal1 s 17070 2054 17106 2395 4 vdd
port 539 nsew
rlabel metal1 s 12078 18145 12114 18486 4 vdd
port 539 nsew
rlabel metal1 s 4590 25255 4626 25596 4 vdd
port 539 nsew
rlabel metal1 s 5838 8665 5874 9006 4 vdd
port 539 nsew
rlabel metal1 s 19086 4715 19122 5056 4 vdd
port 539 nsew
rlabel metal1 s 15822 6295 15858 6636 4 vdd
port 539 nsew
rlabel metal1 s 9102 14694 9138 15035 4 vdd
port 539 nsew
rlabel metal1 s 4590 8665 4626 9006 4 vdd
port 539 nsew
rlabel metal1 s 366 17064 402 17405 4 vdd
port 539 nsew
rlabel metal1 s 846 14985 882 15326 4 vdd
port 539 nsew
rlabel metal1 s 20334 12324 20370 12665 4 vdd
port 539 nsew
rlabel metal1 s 5358 6794 5394 7135 4 vdd
port 539 nsew
rlabel metal1 s 9102 1264 9138 1605 4 vdd
port 539 nsew
rlabel metal1 s 4110 18145 4146 18486 4 vdd
port 539 nsew
rlabel metal1 s 19086 24174 19122 24515 4 vdd
port 539 nsew
rlabel metal1 s 846 9455 882 9796 4 vdd
port 539 nsew
rlabel metal1 s 1614 16274 1650 16615 4 vdd
port 539 nsew
rlabel metal1 s 12078 13904 12114 14245 4 vdd
port 539 nsew
rlabel metal1 s 19566 22095 19602 22436 4 vdd
port 539 nsew
rlabel metal1 s 15822 3634 15858 3975 4 vdd
port 539 nsew
rlabel metal1 s 5838 22885 5874 23226 4 vdd
port 539 nsew
rlabel metal1 s 17838 10744 17874 11085 4 vdd
port 539 nsew
rlabel metal1 s 17070 21804 17106 22145 4 vdd
port 539 nsew
rlabel metal1 s 366 19434 402 19775 4 vdd
port 539 nsew
rlabel metal1 s 18318 11825 18354 12166 4 vdd
port 539 nsew
rlabel metal1 s 1614 5214 1650 5555 4 vdd
port 539 nsew
rlabel metal1 s 3342 5505 3378 5846 4 vdd
port 539 nsew
rlabel metal1 s 3342 13114 3378 13455 4 vdd
port 539 nsew
rlabel metal1 s 7086 23384 7122 23725 4 vdd
port 539 nsew
rlabel metal1 s 13326 13114 13362 13455 4 vdd
port 539 nsew
rlabel metal1 s 20334 1555 20370 1896 4 vdd
port 539 nsew
rlabel metal1 s 12078 20515 12114 20856 4 vdd
port 539 nsew
rlabel metal1 s 7854 18644 7890 18985 4 vdd
port 539 nsew
rlabel metal1 s 19086 5505 19122 5846 4 vdd
port 539 nsew
rlabel metal1 s 17838 7085 17874 7426 4 vdd
port 539 nsew
rlabel metal1 s 16590 18145 16626 18486 4 vdd
port 539 nsew
rlabel metal1 s 7854 11534 7890 11875 4 vdd
port 539 nsew
rlabel metal1 s 7854 9164 7890 9505 4 vdd
port 539 nsew
rlabel metal1 s 9102 16565 9138 16906 4 vdd
port 539 nsew
rlabel metal1 s 11598 4424 11634 4765 4 vdd
port 539 nsew
rlabel metal1 s 2862 2345 2898 2686 4 vdd
port 539 nsew
rlabel metal1 s 2862 474 2898 815 4 vdd
port 539 nsew
rlabel metal1 s 19566 13904 19602 14245 4 vdd
port 539 nsew
rlabel metal1 s 9582 8374 9618 8715 4 vdd
port 539 nsew
rlabel metal1 s 17070 6004 17106 6345 4 vdd
port 539 nsew
rlabel metal1 s 20814 6295 20850 6636 4 vdd
port 539 nsew
rlabel metal1 s 6606 19434 6642 19775 4 vdd
port 539 nsew
rlabel metal1 s 5358 17854 5394 18195 4 vdd
port 539 nsew
rlabel metal1 s 18318 13114 18354 13455 4 vdd
port 539 nsew
rlabel metal1 s 19566 3135 19602 3476 4 vdd
port 539 nsew
rlabel metal1 s 366 18935 402 19276 4 vdd
port 539 nsew
rlabel metal1 s 14574 4715 14610 5056 4 vdd
port 539 nsew
rlabel metal1 s 4590 11825 4626 12166 4 vdd
port 539 nsew
rlabel metal1 s 6606 765 6642 1106 4 vdd
port 539 nsew
rlabel metal1 s 846 21305 882 21646 4 vdd
port 539 nsew
rlabel metal1 s 9102 -25 9138 316 4 vdd
port 539 nsew
rlabel metal1 s 7854 3925 7890 4266 4 vdd
port 539 nsew
rlabel metal1 s 18318 6004 18354 6345 4 vdd
port 539 nsew
rlabel metal1 s 15822 3135 15858 3476 4 vdd
port 539 nsew
rlabel metal1 s 7086 13114 7122 13455 4 vdd
port 539 nsew
rlabel metal1 s 17070 15484 17106 15825 4 vdd
port 539 nsew
rlabel metal1 s 7854 2345 7890 2686 4 vdd
port 539 nsew
rlabel metal1 s 17838 18644 17874 18985 4 vdd
port 539 nsew
rlabel metal1 s 10830 24465 10866 24806 4 vdd
port 539 nsew
rlabel metal1 s 14574 10744 14610 11085 4 vdd
port 539 nsew
rlabel metal1 s 366 2844 402 3185 4 vdd
port 539 nsew
rlabel metal1 s 18318 7584 18354 7925 4 vdd
port 539 nsew
rlabel metal1 s 2094 12615 2130 12956 4 vdd
port 539 nsew
rlabel metal1 s 7086 24465 7122 24806 4 vdd
port 539 nsew
rlabel metal1 s 15822 7875 15858 8216 4 vdd
port 539 nsew
rlabel metal1 s 17070 12615 17106 12956 4 vdd
port 539 nsew
rlabel metal1 s 16590 8665 16626 9006 4 vdd
port 539 nsew
rlabel metal1 s 20814 9164 20850 9505 4 vdd
port 539 nsew
rlabel metal1 s 18318 8665 18354 9006 4 vdd
port 539 nsew
rlabel metal1 s 20814 17355 20850 17696 4 vdd
port 539 nsew
rlabel metal1 s 3342 20515 3378 20856 4 vdd
port 539 nsew
rlabel metal1 s 4590 9455 4626 9796 4 vdd
port 539 nsew
rlabel metal1 s 4110 2844 4146 3185 4 vdd
port 539 nsew
rlabel metal1 s 17070 2844 17106 3185 4 vdd
port 539 nsew
rlabel metal1 s 366 -25 402 316 4 vdd
port 539 nsew
rlabel metal1 s 366 20515 402 20856 4 vdd
port 539 nsew
rlabel metal1 s 8334 22095 8370 22436 4 vdd
port 539 nsew
rlabel metal1 s 17838 19434 17874 19775 4 vdd
port 539 nsew
rlabel metal1 s 15822 5214 15858 5555 4 vdd
port 539 nsew
rlabel metal1 s 6606 11035 6642 11376 4 vdd
port 539 nsew
rlabel metal1 s 19566 11035 19602 11376 4 vdd
port 539 nsew
rlabel metal1 s 4110 5214 4146 5555 4 vdd
port 539 nsew
rlabel metal1 s 18318 1555 18354 1896 4 vdd
port 539 nsew
rlabel metal1 s 14574 2054 14610 2395 4 vdd
port 539 nsew
rlabel metal1 s 15822 23384 15858 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 8374 8370 8715 4 vdd
port 539 nsew
rlabel metal1 s 846 11534 882 11875 4 vdd
port 539 nsew
rlabel metal1 s 16590 6295 16626 6636 4 vdd
port 539 nsew
rlabel metal1 s 5838 24174 5874 24515 4 vdd
port 539 nsew
rlabel metal1 s 12078 6295 12114 6636 4 vdd
port 539 nsew
rlabel metal1 s 846 22885 882 23226 4 vdd
port 539 nsew
rlabel metal1 s 20334 17355 20370 17696 4 vdd
port 539 nsew
rlabel metal1 s 14574 21014 14610 21355 4 vdd
port 539 nsew
rlabel metal1 s 5358 9455 5394 9796 4 vdd
port 539 nsew
rlabel metal1 s 9102 24964 9138 25305 4 vdd
port 539 nsew
rlabel metal1 s 1614 15775 1650 16116 4 vdd
port 539 nsew
rlabel metal1 s 6606 9164 6642 9505 4 vdd
port 539 nsew
rlabel metal1 s 20814 8665 20850 9006 4 vdd
port 539 nsew
rlabel metal1 s 5358 19725 5394 20066 4 vdd
port 539 nsew
rlabel metal1 s 20334 1264 20370 1605 4 vdd
port 539 nsew
rlabel metal1 s 3342 12615 3378 12956 4 vdd
port 539 nsew
rlabel metal1 s 14574 7584 14610 7925 4 vdd
port 539 nsew
rlabel metal1 s 1614 17854 1650 18195 4 vdd
port 539 nsew
rlabel metal1 s 8334 4715 8370 5056 4 vdd
port 539 nsew
rlabel metal1 s 19086 19725 19122 20066 4 vdd
port 539 nsew
rlabel metal1 s 4110 24174 4146 24515 4 vdd
port 539 nsew
rlabel metal1 s 13326 21305 13362 21646 4 vdd
port 539 nsew
rlabel metal1 s 20814 18935 20850 19276 4 vdd
port 539 nsew
rlabel metal1 s 10350 7875 10386 8216 4 vdd
port 539 nsew
rlabel metal1 s 19086 25754 19122 26095 4 vdd
port 539 nsew
rlabel metal1 s 19086 14985 19122 15326 4 vdd
port 539 nsew
rlabel metal1 s 12846 12615 12882 12956 4 vdd
port 539 nsew
rlabel metal1 s 2862 13405 2898 13746 4 vdd
port 539 nsew
rlabel metal1 s 15822 14694 15858 15035 4 vdd
port 539 nsew
rlabel metal1 s 2862 18644 2898 18985 4 vdd
port 539 nsew
rlabel metal1 s 9582 4715 9618 5056 4 vdd
port 539 nsew
rlabel metal1 s 15342 14195 15378 14536 4 vdd
port 539 nsew
rlabel metal1 s 4590 7875 4626 8216 4 vdd
port 539 nsew
rlabel metal1 s 2862 23384 2898 23725 4 vdd
port 539 nsew
rlabel metal1 s 20814 21014 20850 21355 4 vdd
port 539 nsew
rlabel metal1 s 6606 24465 6642 24806 4 vdd
port 539 nsew
rlabel metal1 s 8334 765 8370 1106 4 vdd
port 539 nsew
rlabel metal1 s 9102 20515 9138 20856 4 vdd
port 539 nsew
rlabel metal1 s 19566 1264 19602 1605 4 vdd
port 539 nsew
rlabel metal1 s 9102 12615 9138 12956 4 vdd
port 539 nsew
rlabel metal1 s 4590 3634 4626 3975 4 vdd
port 539 nsew
rlabel metal1 s 3342 25754 3378 26095 4 vdd
port 539 nsew
rlabel metal1 s 366 24174 402 24515 4 vdd
port 539 nsew
rlabel metal1 s 9102 22885 9138 23226 4 vdd
port 539 nsew
rlabel metal1 s 18318 25255 18354 25596 4 vdd
port 539 nsew
rlabel metal1 s 366 8665 402 9006 4 vdd
port 539 nsew
rlabel metal1 s 19086 20515 19122 20856 4 vdd
port 539 nsew
rlabel metal1 s 12846 22594 12882 22935 4 vdd
port 539 nsew
rlabel metal1 s 3342 18935 3378 19276 4 vdd
port 539 nsew
rlabel metal1 s 15342 1264 15378 1605 4 vdd
port 539 nsew
rlabel metal1 s 15342 16565 15378 16906 4 vdd
port 539 nsew
rlabel metal1 s 7854 6295 7890 6636 4 vdd
port 539 nsew
rlabel metal1 s 15342 25754 15378 26095 4 vdd
port 539 nsew
rlabel metal1 s 2094 22594 2130 22935 4 vdd
port 539 nsew
rlabel metal1 s 10350 20224 10386 20565 4 vdd
port 539 nsew
rlabel metal1 s 12846 25255 12882 25596 4 vdd
port 539 nsew
rlabel metal1 s 12846 11035 12882 11376 4 vdd
port 539 nsew
rlabel metal1 s 12846 13405 12882 13746 4 vdd
port 539 nsew
rlabel metal1 s 9102 4715 9138 5056 4 vdd
port 539 nsew
rlabel metal1 s 20814 25754 20850 26095 4 vdd
port 539 nsew
rlabel metal1 s 4590 15775 4626 16116 4 vdd
port 539 nsew
rlabel metal1 s 5838 474 5874 815 4 vdd
port 539 nsew
rlabel metal1 s 19086 17854 19122 18195 4 vdd
port 539 nsew
rlabel metal1 s 15342 5505 15378 5846 4 vdd
port 539 nsew
rlabel metal1 s 10830 14985 10866 15326 4 vdd
port 539 nsew
rlabel metal1 s 2094 6295 2130 6636 4 vdd
port 539 nsew
rlabel metal1 s 17838 9954 17874 10295 4 vdd
port 539 nsew
rlabel metal1 s 12078 19434 12114 19775 4 vdd
port 539 nsew
rlabel metal1 s 19086 14195 19122 14536 4 vdd
port 539 nsew
rlabel metal1 s 1614 7584 1650 7925 4 vdd
port 539 nsew
rlabel metal1 s 16590 5214 16626 5555 4 vdd
port 539 nsew
rlabel metal1 s 7086 12324 7122 12665 4 vdd
port 539 nsew
rlabel metal1 s 9102 11534 9138 11875 4 vdd
port 539 nsew
rlabel metal1 s 366 16565 402 16906 4 vdd
port 539 nsew
rlabel metal1 s 20334 21804 20370 22145 4 vdd
port 539 nsew
rlabel metal1 s 11598 2345 11634 2686 4 vdd
port 539 nsew
rlabel metal1 s 10350 6794 10386 7135 4 vdd
port 539 nsew
rlabel metal1 s 9582 24174 9618 24515 4 vdd
port 539 nsew
rlabel metal1 s 7854 18145 7890 18486 4 vdd
port 539 nsew
rlabel metal1 s 17070 20224 17106 20565 4 vdd
port 539 nsew
rlabel metal1 s 5358 22095 5394 22436 4 vdd
port 539 nsew
rlabel metal1 s 4110 21804 4146 22145 4 vdd
port 539 nsew
rlabel metal1 s 17838 23675 17874 24016 4 vdd
port 539 nsew
rlabel metal1 s 3342 23675 3378 24016 4 vdd
port 539 nsew
rlabel metal1 s 15822 13904 15858 14245 4 vdd
port 539 nsew
rlabel metal1 s 18318 25754 18354 26095 4 vdd
port 539 nsew
rlabel metal1 s 11598 8374 11634 8715 4 vdd
port 539 nsew
rlabel metal1 s 4590 6794 4626 7135 4 vdd
port 539 nsew
rlabel metal1 s 5358 6004 5394 6345 4 vdd
port 539 nsew
rlabel metal1 s 2094 21305 2130 21646 4 vdd
port 539 nsew
rlabel metal1 s 15342 7875 15378 8216 4 vdd
port 539 nsew
rlabel metal1 s 14094 21014 14130 21355 4 vdd
port 539 nsew
rlabel metal1 s 5358 4715 5394 5056 4 vdd
port 539 nsew
rlabel metal1 s 20814 12615 20850 12956 4 vdd
port 539 nsew
rlabel metal1 s 17070 24465 17106 24806 4 vdd
port 539 nsew
rlabel metal1 s 12846 12324 12882 12665 4 vdd
port 539 nsew
rlabel metal1 s 15822 12324 15858 12665 4 vdd
port 539 nsew
rlabel metal1 s 15822 6794 15858 7135 4 vdd
port 539 nsew
rlabel metal1 s 7854 10744 7890 11085 4 vdd
port 539 nsew
rlabel metal1 s 7854 20224 7890 20565 4 vdd
port 539 nsew
rlabel metal1 s 6606 17854 6642 18195 4 vdd
port 539 nsew
rlabel metal1 s 19086 16274 19122 16615 4 vdd
port 539 nsew
rlabel metal1 s 15822 16274 15858 16615 4 vdd
port 539 nsew
rlabel metal1 s 2862 2844 2898 3185 4 vdd
port 539 nsew
rlabel metal1 s 7086 15484 7122 15825 4 vdd
port 539 nsew
rlabel metal1 s 846 20224 882 20565 4 vdd
port 539 nsew
rlabel metal1 s 19086 1555 19122 1896 4 vdd
port 539 nsew
rlabel metal1 s 846 20515 882 20856 4 vdd
port 539 nsew
rlabel metal1 s 10350 17064 10386 17405 4 vdd
port 539 nsew
rlabel metal1 s 846 474 882 815 4 vdd
port 539 nsew
rlabel metal1 s 14094 17854 14130 18195 4 vdd
port 539 nsew
rlabel metal1 s 9102 9455 9138 9796 4 vdd
port 539 nsew
rlabel metal1 s 12846 21804 12882 22145 4 vdd
port 539 nsew
rlabel metal1 s 20334 13904 20370 14245 4 vdd
port 539 nsew
rlabel metal1 s 18318 20515 18354 20856 4 vdd
port 539 nsew
rlabel metal1 s 14574 3135 14610 3476 4 vdd
port 539 nsew
rlabel metal1 s 9582 17854 9618 18195 4 vdd
port 539 nsew
rlabel metal1 s 19086 11035 19122 11376 4 vdd
port 539 nsew
rlabel metal1 s 7854 1264 7890 1605 4 vdd
port 539 nsew
rlabel metal1 s 17838 24465 17874 24806 4 vdd
port 539 nsew
rlabel metal1 s 20334 13114 20370 13455 4 vdd
port 539 nsew
rlabel metal1 s 19566 19725 19602 20066 4 vdd
port 539 nsew
rlabel metal1 s 20334 9164 20370 9505 4 vdd
port 539 nsew
rlabel metal1 s 19566 9455 19602 9796 4 vdd
port 539 nsew
rlabel metal1 s 19566 6794 19602 7135 4 vdd
port 539 nsew
rlabel metal1 s 10830 18935 10866 19276 4 vdd
port 539 nsew
rlabel metal1 s 10350 24964 10386 25305 4 vdd
port 539 nsew
rlabel metal1 s 12078 9164 12114 9505 4 vdd
port 539 nsew
rlabel metal1 s 16590 13114 16626 13455 4 vdd
port 539 nsew
rlabel metal1 s 4590 19725 4626 20066 4 vdd
port 539 nsew
rlabel metal1 s 2094 17355 2130 17696 4 vdd
port 539 nsew
rlabel metal1 s 18318 22095 18354 22436 4 vdd
port 539 nsew
rlabel metal1 s 20814 15484 20850 15825 4 vdd
port 539 nsew
rlabel metal1 s 4590 16274 4626 16615 4 vdd
port 539 nsew
rlabel metal1 s 20814 4424 20850 4765 4 vdd
port 539 nsew
rlabel metal1 s 6606 21305 6642 21646 4 vdd
port 539 nsew
rlabel metal1 s 8334 3925 8370 4266 4 vdd
port 539 nsew
rlabel metal1 s 8334 18145 8370 18486 4 vdd
port 539 nsew
rlabel metal1 s 14574 17355 14610 17696 4 vdd
port 539 nsew
rlabel metal1 s 14094 3634 14130 3975 4 vdd
port 539 nsew
rlabel metal1 s 4110 3135 4146 3476 4 vdd
port 539 nsew
rlabel metal1 s 846 3925 882 4266 4 vdd
port 539 nsew
rlabel metal1 s 17838 6295 17874 6636 4 vdd
port 539 nsew
rlabel metal1 s 9582 5505 9618 5846 4 vdd
port 539 nsew
rlabel metal1 s 14574 18644 14610 18985 4 vdd
port 539 nsew
rlabel metal1 s 3342 7875 3378 8216 4 vdd
port 539 nsew
rlabel metal1 s 14094 2345 14130 2686 4 vdd
port 539 nsew
rlabel metal1 s 846 3634 882 3975 4 vdd
port 539 nsew
rlabel metal1 s 16590 12324 16626 12665 4 vdd
port 539 nsew
rlabel metal1 s 19086 9954 19122 10295 4 vdd
port 539 nsew
rlabel metal1 s 19086 18935 19122 19276 4 vdd
port 539 nsew
rlabel metal1 s 19086 22594 19122 22935 4 vdd
port 539 nsew
rlabel metal1 s 1614 11825 1650 12166 4 vdd
port 539 nsew
rlabel metal1 s 17070 7584 17106 7925 4 vdd
port 539 nsew
rlabel metal1 s 12078 12324 12114 12665 4 vdd
port 539 nsew
rlabel metal1 s 20334 22594 20370 22935 4 vdd
port 539 nsew
rlabel metal1 s 5838 25754 5874 26095 4 vdd
port 539 nsew
rlabel metal1 s 20334 15484 20370 15825 4 vdd
port 539 nsew
rlabel metal1 s 8334 9455 8370 9796 4 vdd
port 539 nsew
rlabel metal1 s 5838 9164 5874 9505 4 vdd
port 539 nsew
rlabel metal1 s 7086 8665 7122 9006 4 vdd
port 539 nsew
rlabel metal1 s 14574 14195 14610 14536 4 vdd
port 539 nsew
rlabel metal1 s 20334 20224 20370 20565 4 vdd
port 539 nsew
rlabel metal1 s 9102 18935 9138 19276 4 vdd
port 539 nsew
rlabel metal1 s 16590 2844 16626 3185 4 vdd
port 539 nsew
rlabel metal1 s 4590 10744 4626 11085 4 vdd
port 539 nsew
rlabel metal1 s 12846 18145 12882 18486 4 vdd
port 539 nsew
rlabel metal1 s 18318 6794 18354 7135 4 vdd
port 539 nsew
rlabel metal1 s 7854 17854 7890 18195 4 vdd
port 539 nsew
rlabel metal1 s 11598 24465 11634 24806 4 vdd
port 539 nsew
rlabel metal1 s 4110 2054 4146 2395 4 vdd
port 539 nsew
rlabel metal1 s 20334 22095 20370 22436 4 vdd
port 539 nsew
rlabel metal1 s 11598 18644 11634 18985 4 vdd
port 539 nsew
rlabel metal1 s 2862 3634 2898 3975 4 vdd
port 539 nsew
rlabel metal1 s 19086 17355 19122 17696 4 vdd
port 539 nsew
rlabel metal1 s 14574 18145 14610 18486 4 vdd
port 539 nsew
rlabel metal1 s 9582 13405 9618 13746 4 vdd
port 539 nsew
rlabel metal1 s 846 18145 882 18486 4 vdd
port 539 nsew
rlabel metal1 s 18318 22885 18354 23226 4 vdd
port 539 nsew
rlabel metal1 s 19086 12324 19122 12665 4 vdd
port 539 nsew
rlabel metal1 s 20334 3634 20370 3975 4 vdd
port 539 nsew
rlabel metal1 s 12078 11035 12114 11376 4 vdd
port 539 nsew
rlabel metal1 s 2862 4715 2898 5056 4 vdd
port 539 nsew
rlabel metal1 s 14094 -25 14130 316 4 vdd
port 539 nsew
rlabel metal1 s 6606 12615 6642 12956 4 vdd
port 539 nsew
rlabel metal1 s 3342 22095 3378 22436 4 vdd
port 539 nsew
rlabel metal1 s 12078 23384 12114 23725 4 vdd
port 539 nsew
rlabel metal1 s 8334 9954 8370 10295 4 vdd
port 539 nsew
rlabel metal1 s 6606 24174 6642 24515 4 vdd
port 539 nsew
rlabel metal1 s 19086 9455 19122 9796 4 vdd
port 539 nsew
rlabel metal1 s 14574 20515 14610 20856 4 vdd
port 539 nsew
rlabel metal1 s 15822 11825 15858 12166 4 vdd
port 539 nsew
rlabel metal1 s 8334 3135 8370 3476 4 vdd
port 539 nsew
rlabel metal1 s 20814 13904 20850 14245 4 vdd
port 539 nsew
rlabel metal1 s 7854 19725 7890 20066 4 vdd
port 539 nsew
rlabel metal1 s 2094 22095 2130 22436 4 vdd
port 539 nsew
rlabel metal1 s 17070 25754 17106 26095 4 vdd
port 539 nsew
rlabel metal1 s 5358 16274 5394 16615 4 vdd
port 539 nsew
rlabel metal1 s 19086 10245 19122 10586 4 vdd
port 539 nsew
rlabel metal1 s 14094 22095 14130 22436 4 vdd
port 539 nsew
rlabel metal1 s 366 5214 402 5555 4 vdd
port 539 nsew
rlabel metal1 s 16590 -25 16626 316 4 vdd
port 539 nsew
rlabel metal1 s 7854 4424 7890 4765 4 vdd
port 539 nsew
rlabel metal1 s 8334 7584 8370 7925 4 vdd
port 539 nsew
rlabel metal1 s 10830 10744 10866 11085 4 vdd
port 539 nsew
rlabel metal1 s 2094 3634 2130 3975 4 vdd
port 539 nsew
rlabel metal1 s 17070 23384 17106 23725 4 vdd
port 539 nsew
rlabel metal1 s 17838 474 17874 815 4 vdd
port 539 nsew
rlabel metal1 s 4110 22594 4146 22935 4 vdd
port 539 nsew
rlabel metal1 s 6606 2345 6642 2686 4 vdd
port 539 nsew
rlabel metal1 s 2094 23675 2130 24016 4 vdd
port 539 nsew
rlabel metal1 s 4110 8374 4146 8715 4 vdd
port 539 nsew
rlabel metal1 s 366 6004 402 6345 4 vdd
port 539 nsew
rlabel metal1 s 4590 24964 4626 25305 4 vdd
port 539 nsew
rlabel metal1 s 16590 7584 16626 7925 4 vdd
port 539 nsew
rlabel metal1 s 19086 12615 19122 12956 4 vdd
port 539 nsew
rlabel metal1 s 19086 1264 19122 1605 4 vdd
port 539 nsew
rlabel metal1 s 2094 15775 2130 16116 4 vdd
port 539 nsew
rlabel metal1 s 16590 3634 16626 3975 4 vdd
port 539 nsew
rlabel metal1 s 5838 12615 5874 12956 4 vdd
port 539 nsew
rlabel metal1 s 8334 13904 8370 14245 4 vdd
port 539 nsew
rlabel metal1 s 9102 19725 9138 20066 4 vdd
port 539 nsew
rlabel metal1 s 4590 11035 4626 11376 4 vdd
port 539 nsew
rlabel metal1 s 2094 1264 2130 1605 4 vdd
port 539 nsew
rlabel metal1 s 17838 17064 17874 17405 4 vdd
port 539 nsew
rlabel metal1 s 366 9164 402 9505 4 vdd
port 539 nsew
rlabel metal1 s 8334 19725 8370 20066 4 vdd
port 539 nsew
rlabel metal1 s 4110 16274 4146 16615 4 vdd
port 539 nsew
rlabel metal1 s 846 9164 882 9505 4 vdd
port 539 nsew
rlabel metal1 s 4110 18935 4146 19276 4 vdd
port 539 nsew
rlabel metal1 s 14574 24174 14610 24515 4 vdd
port 539 nsew
rlabel metal1 s 10830 13405 10866 13746 4 vdd
port 539 nsew
rlabel metal1 s 11598 474 11634 815 4 vdd
port 539 nsew
rlabel metal1 s 10830 9164 10866 9505 4 vdd
port 539 nsew
rlabel metal1 s 17838 23384 17874 23725 4 vdd
port 539 nsew
rlabel metal1 s 1614 19725 1650 20066 4 vdd
port 539 nsew
rlabel metal1 s 846 7875 882 8216 4 vdd
port 539 nsew
rlabel metal1 s 16590 6794 16626 7135 4 vdd
port 539 nsew
rlabel metal1 s 15342 11035 15378 11376 4 vdd
port 539 nsew
rlabel metal1 s 2094 13114 2130 13455 4 vdd
port 539 nsew
rlabel metal1 s 6606 18145 6642 18486 4 vdd
port 539 nsew
rlabel metal1 s 2862 6004 2898 6345 4 vdd
port 539 nsew
rlabel metal1 s 12078 19725 12114 20066 4 vdd
port 539 nsew
rlabel metal1 s 19086 8665 19122 9006 4 vdd
port 539 nsew
rlabel metal1 s 15822 2054 15858 2395 4 vdd
port 539 nsew
rlabel metal1 s 5838 18145 5874 18486 4 vdd
port 539 nsew
rlabel metal1 s 20334 18644 20370 18985 4 vdd
port 539 nsew
rlabel metal1 s 17070 1555 17106 1896 4 vdd
port 539 nsew
rlabel metal1 s 2094 15484 2130 15825 4 vdd
port 539 nsew
rlabel metal1 s 12846 24964 12882 25305 4 vdd
port 539 nsew
rlabel metal1 s 5838 4715 5874 5056 4 vdd
port 539 nsew
rlabel metal1 s 8334 22594 8370 22935 4 vdd
port 539 nsew
rlabel metal1 s 366 24465 402 24806 4 vdd
port 539 nsew
rlabel metal1 s 7854 11825 7890 12166 4 vdd
port 539 nsew
rlabel metal1 s 2094 9164 2130 9505 4 vdd
port 539 nsew
rlabel metal1 s 5358 18644 5394 18985 4 vdd
port 539 nsew
rlabel metal1 s 20814 22885 20850 23226 4 vdd
port 539 nsew
rlabel metal1 s 5358 11534 5394 11875 4 vdd
port 539 nsew
rlabel metal1 s 5358 16565 5394 16906 4 vdd
port 539 nsew
rlabel metal1 s 15822 7584 15858 7925 4 vdd
port 539 nsew
rlabel metal1 s 20814 25255 20850 25596 4 vdd
port 539 nsew
rlabel metal1 s 12078 7584 12114 7925 4 vdd
port 539 nsew
rlabel metal1 s 20814 2345 20850 2686 4 vdd
port 539 nsew
rlabel metal1 s 10350 24465 10386 24806 4 vdd
port 539 nsew
rlabel metal1 s 15342 21305 15378 21646 4 vdd
port 539 nsew
rlabel metal1 s 9102 13405 9138 13746 4 vdd
port 539 nsew
rlabel metal1 s 17838 18145 17874 18486 4 vdd
port 539 nsew
rlabel metal1 s 8334 24964 8370 25305 4 vdd
port 539 nsew
rlabel metal1 s 366 21804 402 22145 4 vdd
port 539 nsew
rlabel metal1 s 14094 21305 14130 21646 4 vdd
port 539 nsew
rlabel metal1 s 7854 25255 7890 25596 4 vdd
port 539 nsew
rlabel metal1 s 846 2345 882 2686 4 vdd
port 539 nsew
rlabel metal1 s 15342 6295 15378 6636 4 vdd
port 539 nsew
rlabel metal1 s 7854 24964 7890 25305 4 vdd
port 539 nsew
rlabel metal1 s 4110 17355 4146 17696 4 vdd
port 539 nsew
rlabel metal1 s 19086 2054 19122 2395 4 vdd
port 539 nsew
rlabel metal1 s 14574 16274 14610 16615 4 vdd
port 539 nsew
rlabel metal1 s 20334 10245 20370 10586 4 vdd
port 539 nsew
rlabel metal1 s 4110 14985 4146 15326 4 vdd
port 539 nsew
rlabel metal1 s 12846 7875 12882 8216 4 vdd
port 539 nsew
rlabel metal1 s 10350 9455 10386 9796 4 vdd
port 539 nsew
rlabel metal1 s 7854 6794 7890 7135 4 vdd
port 539 nsew
rlabel metal1 s 2862 10744 2898 11085 4 vdd
port 539 nsew
rlabel metal1 s 9102 8374 9138 8715 4 vdd
port 539 nsew
rlabel metal1 s 4590 13114 4626 13455 4 vdd
port 539 nsew
rlabel metal1 s 1614 6295 1650 6636 4 vdd
port 539 nsew
rlabel metal1 s 8334 2345 8370 2686 4 vdd
port 539 nsew
rlabel metal1 s 14094 5214 14130 5555 4 vdd
port 539 nsew
rlabel metal1 s 5838 5505 5874 5846 4 vdd
port 539 nsew
rlabel metal1 s 2094 18145 2130 18486 4 vdd
port 539 nsew
rlabel metal1 s 5838 9954 5874 10295 4 vdd
port 539 nsew
rlabel metal1 s 9582 25255 9618 25596 4 vdd
port 539 nsew
rlabel metal1 s 16590 16565 16626 16906 4 vdd
port 539 nsew
rlabel metal1 s 7086 19434 7122 19775 4 vdd
port 539 nsew
rlabel metal1 s 15342 20224 15378 20565 4 vdd
port 539 nsew
rlabel metal1 s 9102 19434 9138 19775 4 vdd
port 539 nsew
rlabel metal1 s 3342 6004 3378 6345 4 vdd
port 539 nsew
rlabel metal1 s 18318 11534 18354 11875 4 vdd
port 539 nsew
rlabel metal1 s 5838 14985 5874 15326 4 vdd
port 539 nsew
rlabel metal1 s 11598 7584 11634 7925 4 vdd
port 539 nsew
rlabel metal1 s 7854 24465 7890 24806 4 vdd
port 539 nsew
rlabel metal1 s 4110 6004 4146 6345 4 vdd
port 539 nsew
rlabel metal1 s 5838 23675 5874 24016 4 vdd
port 539 nsew
rlabel metal1 s 13326 20224 13362 20565 4 vdd
port 539 nsew
rlabel metal1 s 14094 14985 14130 15326 4 vdd
port 539 nsew
rlabel metal1 s 14094 20515 14130 20856 4 vdd
port 539 nsew
rlabel metal1 s 20334 9455 20370 9796 4 vdd
port 539 nsew
rlabel metal1 s 16590 474 16626 815 4 vdd
port 539 nsew
rlabel metal1 s 5358 2054 5394 2395 4 vdd
port 539 nsew
rlabel metal1 s 4110 3925 4146 4266 4 vdd
port 539 nsew
rlabel metal1 s 3342 18145 3378 18486 4 vdd
port 539 nsew
rlabel metal1 s 7854 8665 7890 9006 4 vdd
port 539 nsew
rlabel metal1 s 9582 20515 9618 20856 4 vdd
port 539 nsew
rlabel metal1 s 12846 14195 12882 14536 4 vdd
port 539 nsew
rlabel metal1 s 7854 23384 7890 23725 4 vdd
port 539 nsew
rlabel metal1 s 18318 22594 18354 22935 4 vdd
port 539 nsew
rlabel metal1 s 18318 -25 18354 316 4 vdd
port 539 nsew
rlabel metal1 s 19566 10245 19602 10586 4 vdd
port 539 nsew
rlabel metal1 s 14094 23384 14130 23725 4 vdd
port 539 nsew
rlabel metal1 s 1614 25754 1650 26095 4 vdd
port 539 nsew
rlabel metal1 s 2094 2054 2130 2395 4 vdd
port 539 nsew
rlabel metal1 s 9582 2844 9618 3185 4 vdd
port 539 nsew
rlabel metal1 s 16590 18644 16626 18985 4 vdd
port 539 nsew
rlabel metal1 s 1614 14694 1650 15035 4 vdd
port 539 nsew
rlabel metal1 s 3342 13904 3378 14245 4 vdd
port 539 nsew
rlabel metal1 s 11598 20515 11634 20856 4 vdd
port 539 nsew
rlabel metal1 s 11598 16274 11634 16615 4 vdd
port 539 nsew
rlabel metal1 s 7086 13405 7122 13746 4 vdd
port 539 nsew
rlabel metal1 s 16590 22885 16626 23226 4 vdd
port 539 nsew
rlabel metal1 s 19086 6295 19122 6636 4 vdd
port 539 nsew
rlabel metal1 s 366 25255 402 25596 4 vdd
port 539 nsew
rlabel metal1 s 20814 22594 20850 22935 4 vdd
port 539 nsew
rlabel metal1 s 2094 17854 2130 18195 4 vdd
port 539 nsew
rlabel metal1 s 4590 17355 4626 17696 4 vdd
port 539 nsew
rlabel metal1 s 11598 24174 11634 24515 4 vdd
port 539 nsew
rlabel metal1 s 5358 3634 5394 3975 4 vdd
port 539 nsew
rlabel metal1 s 7854 15484 7890 15825 4 vdd
port 539 nsew
rlabel metal1 s 1614 18935 1650 19276 4 vdd
port 539 nsew
rlabel metal1 s 19086 23384 19122 23725 4 vdd
port 539 nsew
rlabel metal1 s 14574 17854 14610 18195 4 vdd
port 539 nsew
rlabel metal1 s 5358 10245 5394 10586 4 vdd
port 539 nsew
rlabel metal1 s 9582 16565 9618 16906 4 vdd
port 539 nsew
rlabel metal1 s 19086 18145 19122 18486 4 vdd
port 539 nsew
rlabel metal1 s 20814 7085 20850 7426 4 vdd
port 539 nsew
rlabel metal1 s 15822 25255 15858 25596 4 vdd
port 539 nsew
rlabel metal1 s 9582 18935 9618 19276 4 vdd
port 539 nsew
rlabel metal1 s 12078 7875 12114 8216 4 vdd
port 539 nsew
rlabel metal1 s 2094 24465 2130 24806 4 vdd
port 539 nsew
rlabel metal1 s 12846 8665 12882 9006 4 vdd
port 539 nsew
rlabel metal1 s 20814 24964 20850 25305 4 vdd
port 539 nsew
rlabel metal1 s 12846 10744 12882 11085 4 vdd
port 539 nsew
rlabel metal1 s 7854 20515 7890 20856 4 vdd
port 539 nsew
rlabel metal1 s 19086 765 19122 1106 4 vdd
port 539 nsew
rlabel metal1 s 3342 1264 3378 1605 4 vdd
port 539 nsew
rlabel metal1 s 9582 9954 9618 10295 4 vdd
port 539 nsew
rlabel metal1 s 5358 3135 5394 3476 4 vdd
port 539 nsew
rlabel metal1 s 13326 14985 13362 15326 4 vdd
port 539 nsew
rlabel metal1 s 19086 22095 19122 22436 4 vdd
port 539 nsew
rlabel metal1 s 15342 -25 15378 316 4 vdd
port 539 nsew
rlabel metal1 s 6606 13114 6642 13455 4 vdd
port 539 nsew
rlabel metal1 s 8334 20515 8370 20856 4 vdd
port 539 nsew
rlabel metal1 s 1614 11035 1650 11376 4 vdd
port 539 nsew
rlabel metal1 s 2094 5505 2130 5846 4 vdd
port 539 nsew
rlabel metal1 s 366 3135 402 3476 4 vdd
port 539 nsew
rlabel metal1 s 5358 25754 5394 26095 4 vdd
port 539 nsew
rlabel metal1 s 5358 17064 5394 17405 4 vdd
port 539 nsew
rlabel metal1 s 12846 1264 12882 1605 4 vdd
port 539 nsew
rlabel metal1 s 13326 15775 13362 16116 4 vdd
port 539 nsew
rlabel metal1 s 2862 1555 2898 1896 4 vdd
port 539 nsew
rlabel metal1 s 8334 1264 8370 1605 4 vdd
port 539 nsew
rlabel metal1 s 9102 25754 9138 26095 4 vdd
port 539 nsew
rlabel metal1 s 12078 4424 12114 4765 4 vdd
port 539 nsew
rlabel metal1 s 13326 6295 13362 6636 4 vdd
port 539 nsew
rlabel metal1 s 14574 5505 14610 5846 4 vdd
port 539 nsew
rlabel metal1 s 4590 18935 4626 19276 4 vdd
port 539 nsew
rlabel metal1 s 366 18145 402 18486 4 vdd
port 539 nsew
rlabel metal1 s 17838 25754 17874 26095 4 vdd
port 539 nsew
rlabel metal1 s 18318 10245 18354 10586 4 vdd
port 539 nsew
rlabel metal1 s 5838 13114 5874 13455 4 vdd
port 539 nsew
rlabel metal1 s 10350 23675 10386 24016 4 vdd
port 539 nsew
rlabel metal1 s 366 9954 402 10295 4 vdd
port 539 nsew
rlabel metal1 s 14094 20224 14130 20565 4 vdd
port 539 nsew
rlabel metal1 s 10350 8665 10386 9006 4 vdd
port 539 nsew
rlabel metal1 s 9102 17355 9138 17696 4 vdd
port 539 nsew
rlabel metal1 s 20814 12324 20850 12665 4 vdd
port 539 nsew
rlabel metal1 s 4590 22885 4626 23226 4 vdd
port 539 nsew
rlabel metal1 s 16590 9164 16626 9505 4 vdd
port 539 nsew
rlabel metal1 s 7854 2844 7890 3185 4 vdd
port 539 nsew
rlabel metal1 s 2862 9455 2898 9796 4 vdd
port 539 nsew
rlabel metal1 s 15822 2844 15858 3185 4 vdd
port 539 nsew
rlabel metal1 s 6606 1264 6642 1605 4 vdd
port 539 nsew
rlabel metal1 s 10830 5505 10866 5846 4 vdd
port 539 nsew
rlabel metal1 s 10830 2054 10866 2395 4 vdd
port 539 nsew
rlabel metal1 s 2862 24964 2898 25305 4 vdd
port 539 nsew
rlabel metal1 s 18318 2844 18354 3185 4 vdd
port 539 nsew
rlabel metal1 s 3342 18644 3378 18985 4 vdd
port 539 nsew
rlabel metal1 s 8334 13405 8370 13746 4 vdd
port 539 nsew
rlabel metal1 s 3342 23384 3378 23725 4 vdd
port 539 nsew
rlabel metal1 s 10350 16274 10386 16615 4 vdd
port 539 nsew
rlabel metal1 s 6606 11534 6642 11875 4 vdd
port 539 nsew
rlabel metal1 s 1614 4715 1650 5056 4 vdd
port 539 nsew
rlabel metal1 s 2862 20224 2898 20565 4 vdd
port 539 nsew
rlabel metal1 s 9582 25754 9618 26095 4 vdd
port 539 nsew
rlabel metal1 s 20814 2844 20850 3185 4 vdd
port 539 nsew
rlabel metal1 s 19086 7085 19122 7426 4 vdd
port 539 nsew
rlabel metal1 s 5838 1555 5874 1896 4 vdd
port 539 nsew
rlabel metal1 s 12846 5214 12882 5555 4 vdd
port 539 nsew
rlabel metal1 s 11598 7875 11634 8216 4 vdd
port 539 nsew
rlabel metal1 s 12078 765 12114 1106 4 vdd
port 539 nsew
rlabel metal1 s 19566 3925 19602 4266 4 vdd
port 539 nsew
rlabel metal1 s 9102 11035 9138 11376 4 vdd
port 539 nsew
rlabel metal1 s 15822 474 15858 815 4 vdd
port 539 nsew
rlabel metal1 s 12846 4424 12882 4765 4 vdd
port 539 nsew
rlabel metal1 s 11598 9455 11634 9796 4 vdd
port 539 nsew
rlabel metal1 s 4590 4424 4626 4765 4 vdd
port 539 nsew
rlabel metal1 s 15822 13405 15858 13746 4 vdd
port 539 nsew
rlabel metal1 s 14094 474 14130 815 4 vdd
port 539 nsew
rlabel metal1 s 8334 3634 8370 3975 4 vdd
port 539 nsew
rlabel metal1 s 846 8665 882 9006 4 vdd
port 539 nsew
rlabel metal1 s 16590 21305 16626 21646 4 vdd
port 539 nsew
rlabel metal1 s 846 10245 882 10586 4 vdd
port 539 nsew
rlabel metal1 s 20814 1555 20850 1896 4 vdd
port 539 nsew
rlabel metal1 s 15342 2844 15378 3185 4 vdd
port 539 nsew
rlabel metal1 s 15822 1555 15858 1896 4 vdd
port 539 nsew
rlabel metal1 s 19086 6004 19122 6345 4 vdd
port 539 nsew
rlabel metal1 s 17838 1264 17874 1605 4 vdd
port 539 nsew
rlabel metal1 s 17070 12324 17106 12665 4 vdd
port 539 nsew
rlabel metal1 s 846 23675 882 24016 4 vdd
port 539 nsew
rlabel metal1 s 2094 4424 2130 4765 4 vdd
port 539 nsew
rlabel metal1 s 7854 21305 7890 21646 4 vdd
port 539 nsew
rlabel metal1 s 14574 21305 14610 21646 4 vdd
port 539 nsew
rlabel metal1 s 10350 2345 10386 2686 4 vdd
port 539 nsew
rlabel metal1 s 18318 16565 18354 16906 4 vdd
port 539 nsew
rlabel metal2 s 2826 24294 2934 24370 4 gnd
port 541 nsew
rlabel metal2 s 330 5334 438 5410 4 gnd
port 541 nsew
rlabel metal2 s 330 7230 438 7306 4 gnd
port 541 nsew
rlabel metal2 s 10314 21450 10422 21526 4 gnd
port 541 nsew
rlabel metal2 s 330 6914 438 6990 4 gnd
port 541 nsew
rlabel metal2 s 12810 14560 12918 14670 4 gnd
port 541 nsew
rlabel metal2 s 4554 12444 4662 12520 4 gnd
port 541 nsew
rlabel metal2 s 17034 1700 17142 1776 4 gnd
port 541 nsew
rlabel metal2 s 17802 16930 17910 17040 4 gnd
port 541 nsew
rlabel metal2 s 2058 15130 2166 15206 4 gnd
port 541 nsew
rlabel metal2 s 11562 20090 11670 20200 4 gnd
port 541 nsew
rlabel metal2 s 330 14024 438 14100 4 gnd
port 541 nsew
rlabel metal2 s 4074 22460 4182 22570 4 gnd
port 541 nsew
rlabel metal2 s 5322 14340 5430 14416 4 gnd
port 541 nsew
rlabel metal2 s 2058 2174 2166 2250 4 gnd
port 541 nsew
rlabel metal2 s 17802 3280 17910 3356 4 gnd
port 541 nsew
rlabel metal2 s 17802 4860 17910 4936 4 gnd
port 541 nsew
rlabel metal2 s 15306 19554 15414 19630 4 gnd
port 541 nsew
rlabel metal2 s 4074 20344 4182 20420 4 gnd
port 541 nsew
rlabel metal2 s 13290 5080 13398 5190 4 gnd
port 541 nsew
rlabel metal2 s 2826 13550 2934 13626 4 gnd
port 541 nsew
rlabel metal2 s 2058 5650 2166 5726 4 gnd
port 541 nsew
rlabel metal2 s 4074 9284 4182 9360 4 gnd
port 541 nsew
rlabel metal2 s 14538 1384 14646 1460 4 gnd
port 541 nsew
rlabel metal2 s 12810 12444 12918 12520 4 gnd
port 541 nsew
rlabel metal2 s 1578 7230 1686 7306 4 gnd
port 541 nsew
rlabel metal2 s 7050 340 7158 450 4 gnd
port 541 nsew
rlabel metal2 s 10314 16140 10422 16250 4 gnd
port 541 nsew
rlabel metal2 s 5802 15130 5910 15206 4 gnd
port 541 nsew
rlabel metal2 s 17802 15350 17910 15460 4 gnd
port 541 nsew
rlabel metal2 s 11562 1920 11670 2030 4 gnd
port 541 nsew
rlabel metal2 s 2826 20880 2934 20990 4 gnd
port 541 nsew
rlabel metal2 s 6570 9820 6678 9930 4 gnd
port 541 nsew
rlabel metal2 s 17802 25084 17910 25160 4 gnd
port 541 nsew
rlabel metal2 s 7050 17974 7158 18050 4 gnd
port 541 nsew
rlabel metal2 s 11562 12980 11670 13090 4 gnd
port 541 nsew
rlabel metal2 s 7050 24294 7158 24370 4 gnd
port 541 nsew
rlabel metal2 s 4554 11970 4662 12046 4 gnd
port 541 nsew
rlabel metal2 s 19530 20090 19638 20200 4 gnd
port 541 nsew
rlabel metal2 s 2058 7704 2166 7780 4 gnd
port 541 nsew
rlabel metal2 s 14538 10074 14646 10150 4 gnd
port 541 nsew
rlabel metal2 s 4074 21670 4182 21780 4 gnd
port 541 nsew
rlabel metal2 s 7050 15350 7158 15460 4 gnd
port 541 nsew
rlabel metal2 s 20778 15920 20886 15996 4 gnd
port 541 nsew
rlabel metal2 s 15786 9284 15894 9360 4 gnd
port 541 nsew
rlabel metal2 s 8298 10864 8406 10940 4 gnd
port 541 nsew
rlabel metal2 s 15786 12980 15894 13090 4 gnd
port 541 nsew
rlabel metal2 s 10314 12190 10422 12300 4 gnd
port 541 nsew
rlabel metal2 s 7818 12190 7926 12300 4 gnd
port 541 nsew
rlabel metal2 s 7050 9600 7158 9676 4 gnd
port 541 nsew
rlabel metal2 s 15306 25620 15414 25730 4 gnd
port 541 nsew
rlabel metal2 s 330 25620 438 25730 4 gnd
port 541 nsew
rlabel metal2 s 12810 25084 12918 25160 4 gnd
port 541 nsew
rlabel metal2 s 4074 2964 4182 3040 4 gnd
port 541 nsew
rlabel metal2 s 12042 17500 12150 17576 4 gnd
port 541 nsew
rlabel metal2 s 2058 1384 2166 1460 4 gnd
port 541 nsew
rlabel metal2 s 16554 11400 16662 11510 4 gnd
port 541 nsew
rlabel metal2 s 1578 8494 1686 8570 4 gnd
port 541 nsew
rlabel metal2 s 20298 3500 20406 3610 4 gnd
port 541 nsew
rlabel metal2 s 5802 5870 5910 5980 4 gnd
port 541 nsew
rlabel metal2 s 17802 23820 17910 23896 4 gnd
port 541 nsew
rlabel metal2 s 19530 23504 19638 23580 4 gnd
port 541 nsew
rlabel metal2 s 7050 19554 7158 19630 4 gnd
port 541 nsew
rlabel metal2 s 16554 16710 16662 16786 4 gnd
port 541 nsew
rlabel metal2 s 10314 23504 10422 23580 4 gnd
port 541 nsew
rlabel metal2 s 3306 12444 3414 12520 4 gnd
port 541 nsew
rlabel metal2 s 3306 20090 3414 20200 4 gnd
port 541 nsew
rlabel metal2 s 330 11180 438 11256 4 gnd
port 541 nsew
rlabel metal2 s 8298 7230 8406 7306 4 gnd
port 541 nsew
rlabel metal2 s 6570 19870 6678 19946 4 gnd
port 541 nsew
rlabel metal2 s 20298 21134 20406 21210 4 gnd
port 541 nsew
rlabel metal2 s 2058 7230 2166 7306 4 gnd
port 541 nsew
rlabel metal2 s 3306 25874 3414 25950 4 gnd
port 541 nsew
rlabel metal2 s 2058 9030 2166 9140 4 gnd
port 541 nsew
rlabel metal2 s 15786 21134 15894 21210 4 gnd
port 541 nsew
rlabel metal2 s 1578 24610 1686 24686 4 gnd
port 541 nsew
rlabel metal2 s 4554 16710 4662 16786 4 gnd
port 541 nsew
rlabel metal2 s 7050 10390 7158 10466 4 gnd
port 541 nsew
rlabel metal2 s 9066 9030 9174 9140 4 gnd
port 541 nsew
rlabel metal2 s 1578 15920 1686 15996 4 gnd
port 541 nsew
rlabel metal2 s 4074 14560 4182 14670 4 gnd
port 541 nsew
rlabel metal2 s 15306 340 15414 450 4 gnd
port 541 nsew
rlabel metal2 s 15786 15920 15894 15996 4 gnd
port 541 nsew
rlabel metal2 s 20298 25400 20406 25476 4 gnd
port 541 nsew
rlabel metal2 s 11562 9600 11670 9676 4 gnd
port 541 nsew
rlabel metal2 s 19530 13550 19638 13626 4 gnd
port 541 nsew
rlabel metal2 s 17034 4290 17142 4400 4 gnd
port 541 nsew
rlabel metal2 s 7818 15920 7926 15996 4 gnd
port 541 nsew
rlabel metal2 s 12042 9030 12150 9140 4 gnd
port 541 nsew
rlabel metal2 s 19050 4290 19158 4400 4 gnd
port 541 nsew
rlabel metal2 s 6570 24830 6678 24940 4 gnd
port 541 nsew
rlabel metal2 s 330 12444 438 12520 4 gnd
port 541 nsew
rlabel metal2 s 20778 8494 20886 8570 4 gnd
port 541 nsew
rlabel metal2 s 7818 3280 7926 3356 4 gnd
port 541 nsew
rlabel metal2 s 20778 12980 20886 13090 4 gnd
port 541 nsew
rlabel metal2 s 11562 5650 11670 5726 4 gnd
port 541 nsew
rlabel metal2 s 18282 17974 18390 18050 4 gnd
port 541 nsew
rlabel metal2 s 16554 1130 16662 1240 4 gnd
port 541 nsew
rlabel metal2 s 14058 19300 14166 19410 4 gnd
port 541 nsew
rlabel metal2 s 10794 1700 10902 1776 4 gnd
port 541 nsew
rlabel metal2 s 16554 4290 16662 4400 4 gnd
port 541 nsew
rlabel metal2 s 9066 13550 9174 13626 4 gnd
port 541 nsew
rlabel metal2 s 14058 11970 14166 12046 4 gnd
port 541 nsew
rlabel metal2 s 16554 3280 16662 3356 4 gnd
port 541 nsew
rlabel metal2 s 14538 8810 14646 8886 4 gnd
port 541 nsew
rlabel metal2 s 11562 13550 11670 13626 4 gnd
port 541 nsew
rlabel metal2 s 16554 12444 16662 12520 4 gnd
port 541 nsew
rlabel metal2 s 11562 2964 11670 3040 4 gnd
port 541 nsew
rlabel metal2 s 20778 19870 20886 19946 4 gnd
port 541 nsew
rlabel metal2 s 19050 11654 19158 11730 4 gnd
port 541 nsew
rlabel metal2 s 9546 9600 9654 9676 4 gnd
port 541 nsew
rlabel metal2 s 4554 1700 4662 1776 4 gnd
port 541 nsew
rlabel metal2 s 17034 14560 17142 14670 4 gnd
port 541 nsew
rlabel metal2 s 10794 25400 10902 25476 4 gnd
port 541 nsew
rlabel metal2 s 11562 9820 11670 9930 4 gnd
port 541 nsew
rlabel metal2 s 4554 10864 4662 10940 4 gnd
port 541 nsew
rlabel metal2 s 10794 16140 10902 16250 4 gnd
port 541 nsew
rlabel metal2 s 20778 11970 20886 12046 4 gnd
port 541 nsew
rlabel metal2 s 15306 12444 15414 12520 4 gnd
port 541 nsew
rlabel metal2 s 14058 2174 14166 2250 4 gnd
port 541 nsew
rlabel metal2 s 13290 12190 13398 12300 4 gnd
port 541 nsew
rlabel metal2 s 4074 2710 4182 2820 4 gnd
port 541 nsew
rlabel metal2 s 13290 9600 13398 9676 4 gnd
port 541 nsew
rlabel metal2 s 11562 10390 11670 10466 4 gnd
port 541 nsew
rlabel metal2 s 4554 18764 4662 18840 4 gnd
port 541 nsew
rlabel metal2 s 19530 21134 19638 21210 4 gnd
port 541 nsew
rlabel metal2 s 13290 11180 13398 11256 4 gnd
port 541 nsew
rlabel metal2 s 5322 5334 5430 5410 4 gnd
port 541 nsew
rlabel metal2 s 12810 21924 12918 22000 4 gnd
port 541 nsew
rlabel metal2 s 7818 3754 7926 3830 4 gnd
port 541 nsew
rlabel metal2 s 5802 13550 5910 13626 4 gnd
port 541 nsew
rlabel metal2 s 18282 8020 18390 8096 4 gnd
port 541 nsew
rlabel metal2 s 7818 120 7926 196 4 gnd
port 541 nsew
rlabel metal2 s 6570 9284 6678 9360 4 gnd
port 541 nsew
rlabel metal2 s 12810 910 12918 986 4 gnd
port 541 nsew
rlabel metal2 s 9066 15604 9174 15680 4 gnd
port 541 nsew
rlabel metal2 s 19530 23030 19638 23106 4 gnd
port 541 nsew
rlabel metal2 s 7818 22714 7926 22790 4 gnd
port 541 nsew
rlabel metal2 s 7818 25400 7926 25476 4 gnd
port 541 nsew
rlabel metal2 s 18282 10864 18390 10940 4 gnd
port 541 nsew
rlabel metal2 s 7050 1920 7158 2030 4 gnd
port 541 nsew
rlabel metal2 s 15306 6440 15414 6516 4 gnd
port 541 nsew
rlabel metal2 s 4554 22240 4662 22316 4 gnd
port 541 nsew
rlabel metal2 s 4074 1700 4182 1776 4 gnd
port 541 nsew
rlabel metal2 s 9546 3500 9654 3610 4 gnd
port 541 nsew
rlabel metal2 s 810 25620 918 25730 4 gnd
port 541 nsew
rlabel metal2 s 6570 17720 6678 17830 4 gnd
port 541 nsew
rlabel metal2 s 17034 13770 17142 13880 4 gnd
port 541 nsew
rlabel metal2 s 8298 8494 8406 8570 4 gnd
port 541 nsew
rlabel metal2 s 20298 18764 20406 18840 4 gnd
port 541 nsew
rlabel metal2 s 17802 6124 17910 6200 4 gnd
port 541 nsew
rlabel metal2 s 16554 3500 16662 3610 4 gnd
port 541 nsew
rlabel metal2 s 18282 24040 18390 24150 4 gnd
port 541 nsew
rlabel metal2 s 19530 15920 19638 15996 4 gnd
port 541 nsew
rlabel metal2 s 2058 12444 2166 12520 4 gnd
port 541 nsew
rlabel metal2 s 19050 23504 19158 23580 4 gnd
port 541 nsew
rlabel metal2 s 15306 20660 15414 20736 4 gnd
port 541 nsew
rlabel metal2 s 810 8494 918 8570 4 gnd
port 541 nsew
rlabel metal2 s 13290 24610 13398 24686 4 gnd
port 541 nsew
rlabel metal2 s 19530 24610 19638 24686 4 gnd
port 541 nsew
rlabel metal2 s 8298 1384 8406 1460 4 gnd
port 541 nsew
rlabel metal2 s 5322 12190 5430 12300 4 gnd
port 541 nsew
rlabel metal2 s 9546 8240 9654 8350 4 gnd
port 541 nsew
rlabel metal2 s 20778 4290 20886 4400 4 gnd
port 541 nsew
rlabel metal2 s 3306 120 3414 196 4 gnd
port 541 nsew
rlabel metal2 s 330 17500 438 17576 4 gnd
port 541 nsew
rlabel metal2 s 8298 15920 8406 15996 4 gnd
port 541 nsew
rlabel metal2 s 20778 24040 20886 24150 4 gnd
port 541 nsew
rlabel metal2 s 19050 7704 19158 7780 4 gnd
port 541 nsew
rlabel metal2 s 7050 15604 7158 15680 4 gnd
port 541 nsew
rlabel metal2 s 1578 23250 1686 23360 4 gnd
port 541 nsew
rlabel metal2 s 9066 21134 9174 21210 4 gnd
port 541 nsew
rlabel metal2 s 7818 4070 7926 4146 4 gnd
port 541 nsew
rlabel metal2 s 2826 19554 2934 19630 4 gnd
port 541 nsew
rlabel metal2 s 10314 2710 10422 2820 4 gnd
port 541 nsew
rlabel metal2 s 5802 2490 5910 2566 4 gnd
port 541 nsew
rlabel metal2 s 9546 16394 9654 16470 4 gnd
port 541 nsew
rlabel metal2 s 13290 21134 13398 21210 4 gnd
port 541 nsew
rlabel metal2 s 1578 13550 1686 13626 4 gnd
port 541 nsew
rlabel metal2 s 5802 18290 5910 18366 4 gnd
port 541 nsew
rlabel metal2 s 810 14560 918 14670 4 gnd
port 541 nsew
rlabel metal2 s 2058 23030 2166 23106 4 gnd
port 541 nsew
rlabel metal2 s 810 12190 918 12300 4 gnd
port 541 nsew
rlabel metal2 s 7050 120 7158 196 4 gnd
port 541 nsew
rlabel metal2 s 12042 4290 12150 4400 4 gnd
port 541 nsew
rlabel metal2 s 14538 120 14646 196 4 gnd
port 541 nsew
rlabel metal2 s 20778 5650 20886 5726 4 gnd
port 541 nsew
rlabel metal2 s 13290 24830 13398 24940 4 gnd
port 541 nsew
rlabel metal2 s 5802 1130 5910 1240 4 gnd
port 541 nsew
rlabel metal2 s 14538 21450 14646 21526 4 gnd
port 541 nsew
rlabel metal2 s 7818 17974 7926 18050 4 gnd
port 541 nsew
rlabel metal2 s 12042 20344 12150 20420 4 gnd
port 541 nsew
rlabel metal2 s 5802 20880 5910 20990 4 gnd
port 541 nsew
rlabel metal2 s 7050 594 7158 670 4 gnd
port 541 nsew
rlabel metal2 s 17034 4070 17142 4146 4 gnd
port 541 nsew
rlabel metal2 s 18282 20344 18390 20420 4 gnd
port 541 nsew
rlabel metal2 s 15306 3280 15414 3356 4 gnd
port 541 nsew
rlabel metal2 s 10314 17500 10422 17576 4 gnd
port 541 nsew
rlabel metal2 s 10794 3280 10902 3356 4 gnd
port 541 nsew
rlabel metal2 s 5322 6440 5430 6516 4 gnd
port 541 nsew
rlabel metal2 s 10794 23250 10902 23360 4 gnd
port 541 nsew
rlabel metal2 s 19050 9284 19158 9360 4 gnd
port 541 nsew
rlabel metal2 s 14538 6914 14646 6990 4 gnd
port 541 nsew
rlabel metal2 s 330 22714 438 22790 4 gnd
port 541 nsew
rlabel metal2 s 19530 25400 19638 25476 4 gnd
port 541 nsew
rlabel metal2 s 15306 9600 15414 9676 4 gnd
port 541 nsew
rlabel metal2 s 15306 21924 15414 22000 4 gnd
port 541 nsew
rlabel metal2 s 20298 12444 20406 12520 4 gnd
port 541 nsew
rlabel metal2 s 5802 22460 5910 22570 4 gnd
port 541 nsew
rlabel metal2 s 7818 23250 7926 23360 4 gnd
port 541 nsew
rlabel metal2 s 12042 15130 12150 15206 4 gnd
port 541 nsew
rlabel metal2 s 17802 1920 17910 2030 4 gnd
port 541 nsew
rlabel metal2 s 7050 22460 7158 22570 4 gnd
port 541 nsew
rlabel metal2 s 15306 10390 15414 10466 4 gnd
port 541 nsew
rlabel metal2 s 1578 24830 1686 24940 4 gnd
port 541 nsew
rlabel metal2 s 4074 7230 4182 7306 4 gnd
port 541 nsew
rlabel metal2 s 4554 23820 4662 23896 4 gnd
port 541 nsew
rlabel metal2 s 14058 12190 14166 12300 4 gnd
port 541 nsew
rlabel metal2 s 9546 8494 9654 8570 4 gnd
port 541 nsew
rlabel metal2 s 14538 8494 14646 8570 4 gnd
port 541 nsew
rlabel metal2 s 17802 14340 17910 14416 4 gnd
port 541 nsew
rlabel metal2 s 5802 24610 5910 24686 4 gnd
port 541 nsew
rlabel metal2 s 2826 24040 2934 24150 4 gnd
port 541 nsew
rlabel metal2 s 20298 340 20406 450 4 gnd
port 541 nsew
rlabel metal2 s 18282 17184 18390 17260 4 gnd
port 541 nsew
rlabel metal2 s 19530 8494 19638 8570 4 gnd
port 541 nsew
rlabel metal2 s 19050 24294 19158 24370 4 gnd
port 541 nsew
rlabel metal2 s 10314 22460 10422 22570 4 gnd
port 541 nsew
rlabel metal2 s 14538 20344 14646 20420 4 gnd
port 541 nsew
rlabel metal2 s 3306 7704 3414 7780 4 gnd
port 541 nsew
rlabel metal2 s 3306 6914 3414 6990 4 gnd
port 541 nsew
rlabel metal2 s 10314 11180 10422 11256 4 gnd
port 541 nsew
rlabel metal2 s 8298 8240 8406 8350 4 gnd
port 541 nsew
rlabel metal2 s 13290 22460 13398 22570 4 gnd
port 541 nsew
rlabel metal2 s 18282 12444 18390 12520 4 gnd
port 541 nsew
rlabel metal2 s 3306 10864 3414 10940 4 gnd
port 541 nsew
rlabel metal2 s 9066 10390 9174 10466 4 gnd
port 541 nsew
rlabel metal2 s 2058 11400 2166 11510 4 gnd
port 541 nsew
rlabel metal2 s 13290 1384 13398 1460 4 gnd
port 541 nsew
rlabel metal2 s 15786 8240 15894 8350 4 gnd
port 541 nsew
rlabel metal2 s 19530 20344 19638 20420 4 gnd
port 541 nsew
rlabel metal2 s 1578 25400 1686 25476 4 gnd
port 541 nsew
rlabel metal2 s 1578 15604 1686 15680 4 gnd
port 541 nsew
rlabel metal2 s 15306 14340 15414 14416 4 gnd
port 541 nsew
rlabel metal2 s 8298 20344 8406 20420 4 gnd
port 541 nsew
rlabel metal2 s 2826 5870 2934 5980 4 gnd
port 541 nsew
rlabel metal2 s 2826 9284 2934 9360 4 gnd
port 541 nsew
rlabel metal2 s 9546 20660 9654 20736 4 gnd
port 541 nsew
rlabel metal2 s 2826 15920 2934 15996 4 gnd
port 541 nsew
rlabel metal2 s 10794 16710 10902 16786 4 gnd
port 541 nsew
rlabel metal2 s 19530 10390 19638 10466 4 gnd
port 541 nsew
rlabel metal2 s 1578 11180 1686 11256 4 gnd
port 541 nsew
rlabel metal2 s 4554 14340 4662 14416 4 gnd
port 541 nsew
rlabel metal2 s 17034 18290 17142 18366 4 gnd
port 541 nsew
rlabel metal2 s 10794 12190 10902 12300 4 gnd
port 541 nsew
rlabel metal2 s 9066 11970 9174 12046 4 gnd
port 541 nsew
rlabel metal2 s 13290 23820 13398 23896 4 gnd
port 541 nsew
rlabel metal2 s 12042 6914 12150 6990 4 gnd
port 541 nsew
rlabel metal2 s 1578 4290 1686 4400 4 gnd
port 541 nsew
rlabel metal2 s 6570 6124 6678 6200 4 gnd
port 541 nsew
rlabel metal2 s 20298 5650 20406 5726 4 gnd
port 541 nsew
rlabel metal2 s 15786 17184 15894 17260 4 gnd
port 541 nsew
rlabel metal2 s 14058 17500 14166 17576 4 gnd
port 541 nsew
rlabel metal2 s 7050 10074 7158 10150 4 gnd
port 541 nsew
rlabel metal2 s 12810 13234 12918 13310 4 gnd
port 541 nsew
rlabel metal2 s 4554 10610 4662 10720 4 gnd
port 541 nsew
rlabel metal2 s 330 10390 438 10466 4 gnd
port 541 nsew
rlabel metal2 s 17802 14560 17910 14670 4 gnd
port 541 nsew
rlabel metal2 s 810 16930 918 17040 4 gnd
port 541 nsew
rlabel metal2 s 13290 19300 13398 19410 4 gnd
port 541 nsew
rlabel metal2 s 19050 20090 19158 20200 4 gnd
port 541 nsew
rlabel metal2 s 19530 2490 19638 2566 4 gnd
port 541 nsew
rlabel metal2 s 4074 10864 4182 10940 4 gnd
port 541 nsew
rlabel metal2 s 15306 16710 15414 16786 4 gnd
port 541 nsew
rlabel metal2 s 11562 1130 11670 1240 4 gnd
port 541 nsew
rlabel metal2 s 2058 19870 2166 19946 4 gnd
port 541 nsew
rlabel metal2 s 12810 2710 12918 2820 4 gnd
port 541 nsew
rlabel metal2 s 3306 11400 3414 11510 4 gnd
port 541 nsew
rlabel metal2 s 330 3280 438 3356 4 gnd
port 541 nsew
rlabel metal2 s 2058 6660 2166 6770 4 gnd
port 541 nsew
rlabel metal2 s 10314 3500 10422 3610 4 gnd
port 541 nsew
rlabel metal2 s 6570 17500 6678 17576 4 gnd
port 541 nsew
rlabel metal2 s 11562 15130 11670 15206 4 gnd
port 541 nsew
rlabel metal2 s 19530 12190 19638 12300 4 gnd
port 541 nsew
rlabel metal2 s 6570 20660 6678 20736 4 gnd
port 541 nsew
rlabel metal2 s 7050 5870 7158 5980 4 gnd
port 541 nsew
rlabel metal2 s 810 21450 918 21526 4 gnd
port 541 nsew
rlabel metal2 s 11562 22460 11670 22570 4 gnd
port 541 nsew
rlabel metal2 s 1578 9030 1686 9140 4 gnd
port 541 nsew
rlabel metal2 s 15786 13770 15894 13880 4 gnd
port 541 nsew
rlabel metal2 s 330 12980 438 13090 4 gnd
port 541 nsew
rlabel metal2 s 19530 3754 19638 3830 4 gnd
port 541 nsew
rlabel metal2 s 3306 19300 3414 19410 4 gnd
port 541 nsew
rlabel metal2 s 15786 4860 15894 4936 4 gnd
port 541 nsew
rlabel metal2 s 20778 1384 20886 1460 4 gnd
port 541 nsew
rlabel metal2 s 6570 120 6678 196 4 gnd
port 541 nsew
rlabel metal2 s 2058 12760 2166 12836 4 gnd
port 541 nsew
rlabel metal2 s 2058 17720 2166 17830 4 gnd
port 541 nsew
rlabel metal2 s 8298 17974 8406 18050 4 gnd
port 541 nsew
rlabel metal2 s 17802 4070 17910 4146 4 gnd
port 541 nsew
rlabel metal2 s 3306 13770 3414 13880 4 gnd
port 541 nsew
rlabel metal2 s 6570 1920 6678 2030 4 gnd
port 541 nsew
rlabel metal2 s 7818 22240 7926 22316 4 gnd
port 541 nsew
rlabel metal2 s 11562 23504 11670 23580 4 gnd
port 541 nsew
rlabel metal2 s 15306 2490 15414 2566 4 gnd
port 541 nsew
rlabel metal2 s 19530 4290 19638 4400 4 gnd
port 541 nsew
rlabel metal2 s 5322 22240 5430 22316 4 gnd
port 541 nsew
rlabel metal2 s 19530 21450 19638 21526 4 gnd
port 541 nsew
rlabel metal2 s 17034 19080 17142 19156 4 gnd
port 541 nsew
rlabel metal2 s 16554 4860 16662 4936 4 gnd
port 541 nsew
rlabel metal2 s 5802 14814 5910 14890 4 gnd
port 541 nsew
rlabel metal2 s 12042 24610 12150 24686 4 gnd
port 541 nsew
rlabel metal2 s 10314 24294 10422 24370 4 gnd
port 541 nsew
rlabel metal2 s 2826 6124 2934 6200 4 gnd
port 541 nsew
rlabel metal2 s 19530 22460 19638 22570 4 gnd
port 541 nsew
rlabel metal2 s 4074 3754 4182 3830 4 gnd
port 541 nsew
rlabel metal2 s 20298 16140 20406 16250 4 gnd
port 541 nsew
rlabel metal2 s 20298 23820 20406 23896 4 gnd
port 541 nsew
rlabel metal2 s 12810 22240 12918 22316 4 gnd
port 541 nsew
rlabel metal2 s 19530 13770 19638 13880 4 gnd
port 541 nsew
rlabel metal2 s 6570 10610 6678 10720 4 gnd
port 541 nsew
rlabel metal2 s 9546 25620 9654 25730 4 gnd
port 541 nsew
rlabel metal2 s 19530 17184 19638 17260 4 gnd
port 541 nsew
rlabel metal2 s 14538 13770 14646 13880 4 gnd
port 541 nsew
rlabel metal2 s 330 13234 438 13310 4 gnd
port 541 nsew
rlabel metal2 s 10314 15604 10422 15680 4 gnd
port 541 nsew
rlabel metal2 s 10314 14340 10422 14416 4 gnd
port 541 nsew
rlabel metal2 s 5802 21924 5910 22000 4 gnd
port 541 nsew
rlabel metal2 s 7818 24040 7926 24150 4 gnd
port 541 nsew
rlabel metal2 s 12042 19300 12150 19410 4 gnd
port 541 nsew
rlabel metal2 s 330 8240 438 8350 4 gnd
port 541 nsew
rlabel metal2 s 12810 12760 12918 12836 4 gnd
port 541 nsew
rlabel metal2 s 5802 6440 5910 6516 4 gnd
port 541 nsew
rlabel metal2 s 17034 21450 17142 21526 4 gnd
port 541 nsew
rlabel metal2 s 9546 21924 9654 22000 4 gnd
port 541 nsew
rlabel metal2 s 17034 19554 17142 19630 4 gnd
port 541 nsew
rlabel metal2 s 4074 20090 4182 20200 4 gnd
port 541 nsew
rlabel metal2 s 5802 10610 5910 10720 4 gnd
port 541 nsew
rlabel metal2 s 9066 17184 9174 17260 4 gnd
port 541 nsew
rlabel metal2 s 9546 5080 9654 5190 4 gnd
port 541 nsew
rlabel metal2 s 1578 2174 1686 2250 4 gnd
port 541 nsew
rlabel metal2 s 10314 14814 10422 14890 4 gnd
port 541 nsew
rlabel metal2 s 17034 7450 17142 7560 4 gnd
port 541 nsew
rlabel metal2 s 19530 5334 19638 5410 4 gnd
port 541 nsew
rlabel metal2 s 4074 2490 4182 2566 4 gnd
port 541 nsew
rlabel metal2 s 10794 7704 10902 7780 4 gnd
port 541 nsew
rlabel metal2 s 15786 14340 15894 14416 4 gnd
port 541 nsew
rlabel metal2 s 5802 18510 5910 18620 4 gnd
port 541 nsew
rlabel metal2 s 15786 1920 15894 2030 4 gnd
port 541 nsew
rlabel metal2 s 17034 8494 17142 8570 4 gnd
port 541 nsew
rlabel metal2 s 20778 16394 20886 16470 4 gnd
port 541 nsew
rlabel metal2 s 20778 3500 20886 3610 4 gnd
port 541 nsew
rlabel metal2 s 2826 2174 2934 2250 4 gnd
port 541 nsew
rlabel metal2 s 5322 3280 5430 3356 4 gnd
port 541 nsew
rlabel metal2 s 17034 6440 17142 6516 4 gnd
port 541 nsew
rlabel metal2 s 8298 18764 8406 18840 4 gnd
port 541 nsew
rlabel metal2 s 11562 23820 11670 23896 4 gnd
port 541 nsew
rlabel metal2 s 8298 4860 8406 4936 4 gnd
port 541 nsew
rlabel metal2 s 9546 10864 9654 10940 4 gnd
port 541 nsew
rlabel metal2 s 13290 10390 13398 10466 4 gnd
port 541 nsew
rlabel metal2 s 2826 2964 2934 3040 4 gnd
port 541 nsew
rlabel metal2 s 8298 10074 8406 10150 4 gnd
port 541 nsew
rlabel metal2 s 11562 13770 11670 13880 4 gnd
port 541 nsew
rlabel metal2 s 2058 25874 2166 25950 4 gnd
port 541 nsew
rlabel metal2 s 15786 16710 15894 16786 4 gnd
port 541 nsew
rlabel metal2 s 15306 15920 15414 15996 4 gnd
port 541 nsew
rlabel metal2 s 810 14024 918 14100 4 gnd
port 541 nsew
rlabel metal2 s 6570 18764 6678 18840 4 gnd
port 541 nsew
rlabel metal2 s 17034 9820 17142 9930 4 gnd
port 541 nsew
rlabel metal2 s 10314 9600 10422 9676 4 gnd
port 541 nsew
rlabel metal2 s 3306 910 3414 986 4 gnd
port 541 nsew
rlabel metal2 s 4554 13550 4662 13626 4 gnd
port 541 nsew
rlabel metal2 s 8298 594 8406 670 4 gnd
port 541 nsew
rlabel metal2 s 810 2174 918 2250 4 gnd
port 541 nsew
rlabel metal2 s 2826 25084 2934 25160 4 gnd
port 541 nsew
rlabel metal2 s 4074 12980 4182 13090 4 gnd
port 541 nsew
rlabel metal2 s 15306 21450 15414 21526 4 gnd
port 541 nsew
rlabel metal2 s 1578 19554 1686 19630 4 gnd
port 541 nsew
rlabel metal2 s 17802 5650 17910 5726 4 gnd
port 541 nsew
rlabel metal2 s 17034 24830 17142 24940 4 gnd
port 541 nsew
rlabel metal2 s 19530 25084 19638 25160 4 gnd
port 541 nsew
rlabel metal2 s 17034 22240 17142 22316 4 gnd
port 541 nsew
rlabel metal2 s 810 7450 918 7560 4 gnd
port 541 nsew
rlabel metal2 s 14538 5870 14646 5980 4 gnd
port 541 nsew
rlabel metal2 s 7050 2710 7158 2820 4 gnd
port 541 nsew
rlabel metal2 s 20778 19080 20886 19156 4 gnd
port 541 nsew
rlabel metal2 s 5802 7704 5910 7780 4 gnd
port 541 nsew
rlabel metal2 s 17034 12444 17142 12520 4 gnd
port 541 nsew
rlabel metal2 s 15786 8020 15894 8096 4 gnd
port 541 nsew
rlabel metal2 s 14058 3280 14166 3356 4 gnd
port 541 nsew
rlabel metal2 s 12042 5080 12150 5190 4 gnd
port 541 nsew
rlabel metal2 s 20298 24830 20406 24940 4 gnd
port 541 nsew
rlabel metal2 s 5802 11180 5910 11256 4 gnd
port 541 nsew
rlabel metal2 s 16554 8240 16662 8350 4 gnd
port 541 nsew
rlabel metal2 s 20298 2174 20406 2250 4 gnd
port 541 nsew
rlabel metal2 s 4074 14814 4182 14890 4 gnd
port 541 nsew
rlabel metal2 s 18282 7230 18390 7306 4 gnd
port 541 nsew
rlabel metal2 s 20298 15604 20406 15680 4 gnd
port 541 nsew
rlabel metal2 s 9066 14024 9174 14100 4 gnd
port 541 nsew
rlabel metal2 s 9546 1130 9654 1240 4 gnd
port 541 nsew
rlabel metal2 s 9546 13550 9654 13626 4 gnd
port 541 nsew
rlabel metal2 s 20778 12760 20886 12836 4 gnd
port 541 nsew
rlabel metal2 s 330 17974 438 18050 4 gnd
port 541 nsew
rlabel metal2 s 14058 19870 14166 19946 4 gnd
port 541 nsew
rlabel metal2 s 18282 3280 18390 3356 4 gnd
port 541 nsew
rlabel metal2 s 16554 18764 16662 18840 4 gnd
port 541 nsew
rlabel metal2 s 12810 20090 12918 20200 4 gnd
port 541 nsew
rlabel metal2 s 7818 1130 7926 1240 4 gnd
port 541 nsew
rlabel metal2 s 19530 16394 19638 16470 4 gnd
port 541 nsew
rlabel metal2 s 7818 16394 7926 16470 4 gnd
port 541 nsew
rlabel metal2 s 17034 5080 17142 5190 4 gnd
port 541 nsew
rlabel metal2 s 3306 16710 3414 16786 4 gnd
port 541 nsew
rlabel metal2 s 6570 910 6678 986 4 gnd
port 541 nsew
rlabel metal2 s 20298 14560 20406 14670 4 gnd
port 541 nsew
rlabel metal2 s 11562 6124 11670 6200 4 gnd
port 541 nsew
rlabel metal2 s 19530 2710 19638 2820 4 gnd
port 541 nsew
rlabel metal2 s 15786 6124 15894 6200 4 gnd
port 541 nsew
rlabel metal2 s 5322 12760 5430 12836 4 gnd
port 541 nsew
rlabel metal2 s 17802 19080 17910 19156 4 gnd
port 541 nsew
rlabel metal2 s 20298 25084 20406 25160 4 gnd
port 541 nsew
rlabel metal2 s 3306 9600 3414 9676 4 gnd
port 541 nsew
rlabel metal2 s 11562 13234 11670 13310 4 gnd
port 541 nsew
rlabel metal2 s 2058 25620 2166 25730 4 gnd
port 541 nsew
rlabel metal2 s 19050 18510 19158 18620 4 gnd
port 541 nsew
rlabel metal2 s 20298 5870 20406 5980 4 gnd
port 541 nsew
rlabel metal2 s 18282 20090 18390 20200 4 gnd
port 541 nsew
rlabel metal2 s 14058 10610 14166 10720 4 gnd
port 541 nsew
rlabel metal2 s 4074 1130 4182 1240 4 gnd
port 541 nsew
rlabel metal2 s 17034 22714 17142 22790 4 gnd
port 541 nsew
rlabel metal2 s 5322 16930 5430 17040 4 gnd
port 541 nsew
rlabel metal2 s 5322 6124 5430 6200 4 gnd
port 541 nsew
rlabel metal2 s 15306 4070 15414 4146 4 gnd
port 541 nsew
rlabel metal2 s 2058 17974 2166 18050 4 gnd
port 541 nsew
rlabel metal2 s 3306 1700 3414 1776 4 gnd
port 541 nsew
rlabel metal2 s 20778 6440 20886 6516 4 gnd
port 541 nsew
rlabel metal2 s 2058 120 2166 196 4 gnd
port 541 nsew
rlabel metal2 s 19530 7704 19638 7780 4 gnd
port 541 nsew
rlabel metal2 s 17802 19300 17910 19410 4 gnd
port 541 nsew
rlabel metal2 s 15306 15604 15414 15680 4 gnd
port 541 nsew
rlabel metal2 s 8298 5334 8406 5410 4 gnd
port 541 nsew
rlabel metal2 s 15306 17184 15414 17260 4 gnd
port 541 nsew
rlabel metal2 s 7818 1700 7926 1776 4 gnd
port 541 nsew
rlabel metal2 s 19530 15130 19638 15206 4 gnd
port 541 nsew
rlabel metal2 s 12810 14024 12918 14100 4 gnd
port 541 nsew
rlabel metal2 s 15306 14024 15414 14100 4 gnd
port 541 nsew
rlabel metal2 s 7818 22460 7926 22570 4 gnd
port 541 nsew
rlabel metal2 s 10794 14560 10902 14670 4 gnd
port 541 nsew
rlabel metal2 s 17802 12760 17910 12836 4 gnd
port 541 nsew
rlabel metal2 s 4554 11180 4662 11256 4 gnd
port 541 nsew
rlabel metal2 s 7818 8240 7926 8350 4 gnd
port 541 nsew
rlabel metal2 s 10314 15350 10422 15460 4 gnd
port 541 nsew
rlabel metal2 s 10314 594 10422 670 4 gnd
port 541 nsew
rlabel metal2 s 17802 12444 17910 12520 4 gnd
port 541 nsew
rlabel metal2 s 12810 6914 12918 6990 4 gnd
port 541 nsew
rlabel metal2 s 20298 22460 20406 22570 4 gnd
port 541 nsew
rlabel metal2 s 12810 25400 12918 25476 4 gnd
port 541 nsew
rlabel metal2 s 14538 16140 14646 16250 4 gnd
port 541 nsew
rlabel metal2 s 4554 11654 4662 11730 4 gnd
port 541 nsew
rlabel metal2 s 2058 10390 2166 10466 4 gnd
port 541 nsew
rlabel metal2 s 15786 23504 15894 23580 4 gnd
port 541 nsew
rlabel metal2 s 1578 2490 1686 2566 4 gnd
port 541 nsew
rlabel metal2 s 18282 4070 18390 4146 4 gnd
port 541 nsew
rlabel metal2 s 17034 4544 17142 4620 4 gnd
port 541 nsew
rlabel metal2 s 10794 11400 10902 11510 4 gnd
port 541 nsew
rlabel metal2 s 14058 17974 14166 18050 4 gnd
port 541 nsew
rlabel metal2 s 12042 14024 12150 14100 4 gnd
port 541 nsew
rlabel metal2 s 17802 10610 17910 10720 4 gnd
port 541 nsew
rlabel metal2 s 19050 2490 19158 2566 4 gnd
port 541 nsew
rlabel metal2 s 810 11400 918 11510 4 gnd
port 541 nsew
rlabel metal2 s 9546 19300 9654 19410 4 gnd
port 541 nsew
rlabel metal2 s 2058 24610 2166 24686 4 gnd
port 541 nsew
rlabel metal2 s 4074 18290 4182 18366 4 gnd
port 541 nsew
rlabel metal2 s 9546 5650 9654 5726 4 gnd
port 541 nsew
rlabel metal2 s 6570 14340 6678 14416 4 gnd
port 541 nsew
rlabel metal2 s 2058 15920 2166 15996 4 gnd
port 541 nsew
rlabel metal2 s 9066 4860 9174 4936 4 gnd
port 541 nsew
rlabel metal2 s 810 14340 918 14416 4 gnd
port 541 nsew
rlabel metal2 s 2058 14340 2166 14416 4 gnd
port 541 nsew
rlabel metal2 s 7818 10610 7926 10720 4 gnd
port 541 nsew
rlabel metal2 s 14538 16930 14646 17040 4 gnd
port 541 nsew
rlabel metal2 s 330 25874 438 25950 4 gnd
port 541 nsew
rlabel metal2 s 6570 7230 6678 7306 4 gnd
port 541 nsew
rlabel metal2 s 3306 24040 3414 24150 4 gnd
port 541 nsew
rlabel metal2 s 2826 16140 2934 16250 4 gnd
port 541 nsew
rlabel metal2 s 11562 14814 11670 14890 4 gnd
port 541 nsew
rlabel metal2 s 10314 1700 10422 1776 4 gnd
port 541 nsew
rlabel metal2 s 5802 4860 5910 4936 4 gnd
port 541 nsew
rlabel metal2 s 18282 9284 18390 9360 4 gnd
port 541 nsew
rlabel metal2 s 2826 11970 2934 12046 4 gnd
port 541 nsew
rlabel metal2 s 14538 24830 14646 24940 4 gnd
port 541 nsew
rlabel metal2 s 10794 14814 10902 14890 4 gnd
port 541 nsew
rlabel metal2 s 19530 11180 19638 11256 4 gnd
port 541 nsew
rlabel metal2 s 3306 25620 3414 25730 4 gnd
port 541 nsew
rlabel metal2 s 16554 120 16662 196 4 gnd
port 541 nsew
rlabel metal2 s 15306 5870 15414 5980 4 gnd
port 541 nsew
rlabel metal2 s 2826 9820 2934 9930 4 gnd
port 541 nsew
rlabel metal2 s 5802 6660 5910 6770 4 gnd
port 541 nsew
rlabel metal2 s 9066 5080 9174 5190 4 gnd
port 541 nsew
rlabel metal2 s 810 17720 918 17830 4 gnd
port 541 nsew
rlabel metal2 s 3306 20880 3414 20990 4 gnd
port 541 nsew
rlabel metal2 s 2826 25620 2934 25730 4 gnd
port 541 nsew
rlabel metal2 s 10794 2964 10902 3040 4 gnd
port 541 nsew
rlabel metal2 s 1578 17974 1686 18050 4 gnd
port 541 nsew
rlabel metal2 s 2058 24294 2166 24370 4 gnd
port 541 nsew
rlabel metal2 s 4074 24294 4182 24370 4 gnd
port 541 nsew
rlabel metal2 s 20298 15130 20406 15206 4 gnd
port 541 nsew
rlabel metal2 s 13290 1130 13398 1240 4 gnd
port 541 nsew
rlabel metal2 s 15786 4290 15894 4400 4 gnd
port 541 nsew
rlabel metal2 s 7050 23820 7158 23896 4 gnd
port 541 nsew
rlabel metal2 s 12810 1920 12918 2030 4 gnd
port 541 nsew
rlabel metal2 s 7818 2174 7926 2250 4 gnd
port 541 nsew
rlabel metal2 s 12042 1700 12150 1776 4 gnd
port 541 nsew
rlabel metal2 s 12042 10074 12150 10150 4 gnd
port 541 nsew
rlabel metal2 s 20298 14024 20406 14100 4 gnd
port 541 nsew
rlabel metal2 s 5802 2710 5910 2820 4 gnd
port 541 nsew
rlabel metal2 s 19530 12980 19638 13090 4 gnd
port 541 nsew
rlabel metal2 s 11562 19870 11670 19946 4 gnd
port 541 nsew
rlabel metal2 s 14538 9600 14646 9676 4 gnd
port 541 nsew
rlabel metal2 s 9066 10864 9174 10940 4 gnd
port 541 nsew
rlabel metal2 s 12810 6440 12918 6516 4 gnd
port 541 nsew
rlabel metal2 s 14538 10390 14646 10466 4 gnd
port 541 nsew
rlabel metal2 s 9546 2710 9654 2820 4 gnd
port 541 nsew
rlabel metal2 s 14058 23504 14166 23580 4 gnd
port 541 nsew
rlabel metal2 s 17034 12760 17142 12836 4 gnd
port 541 nsew
rlabel metal2 s 15306 23820 15414 23896 4 gnd
port 541 nsew
rlabel metal2 s 20778 6124 20886 6200 4 gnd
port 541 nsew
rlabel metal2 s 11562 9284 11670 9360 4 gnd
port 541 nsew
rlabel metal2 s 14538 5650 14646 5726 4 gnd
port 541 nsew
rlabel metal2 s 5322 8240 5430 8350 4 gnd
port 541 nsew
rlabel metal2 s 16554 25084 16662 25160 4 gnd
port 541 nsew
rlabel metal2 s 17802 8810 17910 8886 4 gnd
port 541 nsew
rlabel metal2 s 10314 9284 10422 9360 4 gnd
port 541 nsew
rlabel metal2 s 20298 20880 20406 20990 4 gnd
port 541 nsew
rlabel metal2 s 10314 16710 10422 16786 4 gnd
port 541 nsew
rlabel metal2 s 15786 910 15894 986 4 gnd
port 541 nsew
rlabel metal2 s 5802 16140 5910 16250 4 gnd
port 541 nsew
rlabel metal2 s 14538 22460 14646 22570 4 gnd
port 541 nsew
rlabel metal2 s 17802 6440 17910 6516 4 gnd
port 541 nsew
rlabel metal2 s 7050 19870 7158 19946 4 gnd
port 541 nsew
rlabel metal2 s 18282 3500 18390 3610 4 gnd
port 541 nsew
rlabel metal2 s 15306 13234 15414 13310 4 gnd
port 541 nsew
rlabel metal2 s 7050 17500 7158 17576 4 gnd
port 541 nsew
rlabel metal2 s 11562 19080 11670 19156 4 gnd
port 541 nsew
rlabel metal2 s 330 6660 438 6770 4 gnd
port 541 nsew
rlabel metal2 s 20778 7450 20886 7560 4 gnd
port 541 nsew
rlabel metal2 s 14538 19554 14646 19630 4 gnd
port 541 nsew
rlabel metal2 s 20778 4070 20886 4146 4 gnd
port 541 nsew
rlabel metal2 s 5322 7450 5430 7560 4 gnd
port 541 nsew
rlabel metal2 s 16554 15130 16662 15206 4 gnd
port 541 nsew
rlabel metal2 s 14538 7450 14646 7560 4 gnd
port 541 nsew
rlabel metal2 s 15786 13234 15894 13310 4 gnd
port 541 nsew
rlabel metal2 s 330 120 438 196 4 gnd
port 541 nsew
rlabel metal2 s 17034 25874 17142 25950 4 gnd
port 541 nsew
rlabel metal2 s 9066 3500 9174 3610 4 gnd
port 541 nsew
rlabel metal2 s 20298 2964 20406 3040 4 gnd
port 541 nsew
rlabel metal2 s 10314 2490 10422 2566 4 gnd
port 541 nsew
rlabel metal2 s 3306 8240 3414 8350 4 gnd
port 541 nsew
rlabel metal2 s 20298 1920 20406 2030 4 gnd
port 541 nsew
rlabel metal2 s 17802 9820 17910 9930 4 gnd
port 541 nsew
rlabel metal2 s 7050 10864 7158 10940 4 gnd
port 541 nsew
rlabel metal2 s 2826 12190 2934 12300 4 gnd
port 541 nsew
rlabel metal2 s 810 10074 918 10150 4 gnd
port 541 nsew
rlabel metal2 s 18282 12980 18390 13090 4 gnd
port 541 nsew
rlabel metal2 s 4074 17184 4182 17260 4 gnd
port 541 nsew
rlabel metal2 s 2826 1384 2934 1460 4 gnd
port 541 nsew
rlabel metal2 s 18282 120 18390 196 4 gnd
port 541 nsew
rlabel metal2 s 7818 20880 7926 20990 4 gnd
port 541 nsew
rlabel metal2 s 16554 340 16662 450 4 gnd
port 541 nsew
rlabel metal2 s 330 19080 438 19156 4 gnd
port 541 nsew
rlabel metal2 s 18282 8810 18390 8886 4 gnd
port 541 nsew
rlabel metal2 s 810 9284 918 9360 4 gnd
port 541 nsew
rlabel metal2 s 5802 23820 5910 23896 4 gnd
port 541 nsew
rlabel metal2 s 3306 18290 3414 18366 4 gnd
port 541 nsew
rlabel metal2 s 18282 10390 18390 10466 4 gnd
port 541 nsew
rlabel metal2 s 3306 17500 3414 17576 4 gnd
port 541 nsew
rlabel metal2 s 5322 14560 5430 14670 4 gnd
port 541 nsew
rlabel metal2 s 20778 18510 20886 18620 4 gnd
port 541 nsew
rlabel metal2 s 810 25874 918 25950 4 gnd
port 541 nsew
rlabel metal2 s 19530 14340 19638 14416 4 gnd
port 541 nsew
rlabel metal2 s 5802 13234 5910 13310 4 gnd
port 541 nsew
rlabel metal2 s 4074 13770 4182 13880 4 gnd
port 541 nsew
rlabel metal2 s 9066 19870 9174 19946 4 gnd
port 541 nsew
rlabel metal2 s 16554 19554 16662 19630 4 gnd
port 541 nsew
rlabel metal2 s 5322 16394 5430 16470 4 gnd
port 541 nsew
rlabel metal2 s 14058 21450 14166 21526 4 gnd
port 541 nsew
rlabel metal2 s 12810 18290 12918 18366 4 gnd
port 541 nsew
rlabel metal2 s 5802 5080 5910 5190 4 gnd
port 541 nsew
rlabel metal2 s 810 1700 918 1776 4 gnd
port 541 nsew
rlabel metal2 s 810 19554 918 19630 4 gnd
port 541 nsew
rlabel metal2 s 11562 6914 11670 6990 4 gnd
port 541 nsew
rlabel metal2 s 14058 20344 14166 20420 4 gnd
port 541 nsew
rlabel metal2 s 5322 24040 5430 24150 4 gnd
port 541 nsew
rlabel metal2 s 12810 16140 12918 16250 4 gnd
port 541 nsew
rlabel metal2 s 7818 7230 7926 7306 4 gnd
port 541 nsew
rlabel metal2 s 13290 25874 13398 25950 4 gnd
port 541 nsew
rlabel metal2 s 2826 8240 2934 8350 4 gnd
port 541 nsew
rlabel metal2 s 17034 14340 17142 14416 4 gnd
port 541 nsew
rlabel metal2 s 4554 8020 4662 8096 4 gnd
port 541 nsew
rlabel metal2 s 7050 24610 7158 24686 4 gnd
port 541 nsew
rlabel metal2 s 19050 19300 19158 19410 4 gnd
port 541 nsew
rlabel metal2 s 2826 594 2934 670 4 gnd
port 541 nsew
rlabel metal2 s 9546 8810 9654 8886 4 gnd
port 541 nsew
rlabel metal2 s 18282 23030 18390 23106 4 gnd
port 541 nsew
rlabel metal2 s 11562 25084 11670 25160 4 gnd
port 541 nsew
rlabel metal2 s 17802 5870 17910 5980 4 gnd
port 541 nsew
rlabel metal2 s 15306 24294 15414 24370 4 gnd
port 541 nsew
rlabel metal2 s 10314 14024 10422 14100 4 gnd
port 541 nsew
rlabel metal2 s 19050 10390 19158 10466 4 gnd
port 541 nsew
rlabel metal2 s 11562 17974 11670 18050 4 gnd
port 541 nsew
rlabel metal2 s 330 10074 438 10150 4 gnd
port 541 nsew
rlabel metal2 s 16554 13770 16662 13880 4 gnd
port 541 nsew
rlabel metal2 s 20778 25874 20886 25950 4 gnd
port 541 nsew
rlabel metal2 s 7050 18764 7158 18840 4 gnd
port 541 nsew
rlabel metal2 s 2058 25400 2166 25476 4 gnd
port 541 nsew
rlabel metal2 s 11562 24040 11670 24150 4 gnd
port 541 nsew
rlabel metal2 s 8298 12190 8406 12300 4 gnd
port 541 nsew
rlabel metal2 s 19530 17974 19638 18050 4 gnd
port 541 nsew
rlabel metal2 s 11562 8240 11670 8350 4 gnd
port 541 nsew
rlabel metal2 s 330 22460 438 22570 4 gnd
port 541 nsew
rlabel metal2 s 15306 10610 15414 10720 4 gnd
port 541 nsew
rlabel metal2 s 17802 8494 17910 8570 4 gnd
port 541 nsew
rlabel metal2 s 20778 12190 20886 12300 4 gnd
port 541 nsew
rlabel metal2 s 4554 17974 4662 18050 4 gnd
port 541 nsew
rlabel metal2 s 9546 6914 9654 6990 4 gnd
port 541 nsew
rlabel metal2 s 15786 20880 15894 20990 4 gnd
port 541 nsew
rlabel metal2 s 12042 2490 12150 2566 4 gnd
port 541 nsew
rlabel metal2 s 14058 14814 14166 14890 4 gnd
port 541 nsew
rlabel metal2 s 13290 8020 13398 8096 4 gnd
port 541 nsew
rlabel metal2 s 5802 340 5910 450 4 gnd
port 541 nsew
rlabel metal2 s 8298 16140 8406 16250 4 gnd
port 541 nsew
rlabel metal2 s 19530 11970 19638 12046 4 gnd
port 541 nsew
rlabel metal2 s 20298 6440 20406 6516 4 gnd
port 541 nsew
rlabel metal2 s 4554 1384 4662 1460 4 gnd
port 541 nsew
rlabel metal2 s 18282 6440 18390 6516 4 gnd
port 541 nsew
rlabel metal2 s 2826 11654 2934 11730 4 gnd
port 541 nsew
rlabel metal2 s 20298 8494 20406 8570 4 gnd
port 541 nsew
rlabel metal2 s 7050 11180 7158 11256 4 gnd
port 541 nsew
rlabel metal2 s 5322 14814 5430 14890 4 gnd
port 541 nsew
rlabel metal2 s 810 20344 918 20420 4 gnd
port 541 nsew
rlabel metal2 s 5322 12444 5430 12520 4 gnd
port 541 nsew
rlabel metal2 s 20298 23250 20406 23360 4 gnd
port 541 nsew
rlabel metal2 s 330 1130 438 1240 4 gnd
port 541 nsew
rlabel metal2 s 14058 23030 14166 23106 4 gnd
port 541 nsew
rlabel metal2 s 5802 22714 5910 22790 4 gnd
port 541 nsew
rlabel metal2 s 20298 16394 20406 16470 4 gnd
port 541 nsew
rlabel metal2 s 10794 4070 10902 4146 4 gnd
port 541 nsew
rlabel metal2 s 14538 8020 14646 8096 4 gnd
port 541 nsew
rlabel metal2 s 17034 7230 17142 7306 4 gnd
port 541 nsew
rlabel metal2 s 15786 22460 15894 22570 4 gnd
port 541 nsew
rlabel metal2 s 13290 8240 13398 8350 4 gnd
port 541 nsew
rlabel metal2 s 11562 24610 11670 24686 4 gnd
port 541 nsew
rlabel metal2 s 5802 11970 5910 12046 4 gnd
port 541 nsew
rlabel metal2 s 810 20090 918 20200 4 gnd
port 541 nsew
rlabel metal2 s 13290 4290 13398 4400 4 gnd
port 541 nsew
rlabel metal2 s 3306 11970 3414 12046 4 gnd
port 541 nsew
rlabel metal2 s 5802 23030 5910 23106 4 gnd
port 541 nsew
rlabel metal2 s 20298 21924 20406 22000 4 gnd
port 541 nsew
rlabel metal2 s 2058 11970 2166 12046 4 gnd
port 541 nsew
rlabel metal2 s 15786 24040 15894 24150 4 gnd
port 541 nsew
rlabel metal2 s 10314 17974 10422 18050 4 gnd
port 541 nsew
rlabel metal2 s 13290 3500 13398 3610 4 gnd
port 541 nsew
rlabel metal2 s 18282 15604 18390 15680 4 gnd
port 541 nsew
rlabel metal2 s 7818 11970 7926 12046 4 gnd
port 541 nsew
rlabel metal2 s 8298 18510 8406 18620 4 gnd
port 541 nsew
rlabel metal2 s 4074 3500 4182 3610 4 gnd
port 541 nsew
rlabel metal2 s 19050 25874 19158 25950 4 gnd
port 541 nsew
rlabel metal2 s 7050 1700 7158 1776 4 gnd
port 541 nsew
rlabel metal2 s 14058 12760 14166 12836 4 gnd
port 541 nsew
rlabel metal2 s 18282 9600 18390 9676 4 gnd
port 541 nsew
rlabel metal2 s 15306 8020 15414 8096 4 gnd
port 541 nsew
rlabel metal2 s 18282 23820 18390 23896 4 gnd
port 541 nsew
rlabel metal2 s 10794 8810 10902 8886 4 gnd
port 541 nsew
rlabel metal2 s 19050 1130 19158 1240 4 gnd
port 541 nsew
rlabel metal2 s 14058 9030 14166 9140 4 gnd
port 541 nsew
rlabel metal2 s 15306 18510 15414 18620 4 gnd
port 541 nsew
rlabel metal2 s 810 7704 918 7780 4 gnd
port 541 nsew
rlabel metal2 s 5322 19554 5430 19630 4 gnd
port 541 nsew
rlabel metal2 s 8298 21924 8406 22000 4 gnd
port 541 nsew
rlabel metal2 s 19050 16930 19158 17040 4 gnd
port 541 nsew
rlabel metal2 s 20778 120 20886 196 4 gnd
port 541 nsew
rlabel metal2 s 17034 16930 17142 17040 4 gnd
port 541 nsew
rlabel metal2 s 10794 18290 10902 18366 4 gnd
port 541 nsew
rlabel metal2 s 19530 23820 19638 23896 4 gnd
port 541 nsew
rlabel metal2 s 4074 4070 4182 4146 4 gnd
port 541 nsew
rlabel metal2 s 12810 23504 12918 23580 4 gnd
port 541 nsew
rlabel metal2 s 9546 1700 9654 1776 4 gnd
port 541 nsew
rlabel metal2 s 12810 21134 12918 21210 4 gnd
port 541 nsew
rlabel metal2 s 7818 7704 7926 7780 4 gnd
port 541 nsew
rlabel metal2 s 8298 12444 8406 12520 4 gnd
port 541 nsew
rlabel metal2 s 10794 13234 10902 13310 4 gnd
port 541 nsew
rlabel metal2 s 7818 9600 7926 9676 4 gnd
port 541 nsew
rlabel metal2 s 16554 6914 16662 6990 4 gnd
port 541 nsew
rlabel metal2 s 12810 10864 12918 10940 4 gnd
port 541 nsew
rlabel metal2 s 7818 14340 7926 14416 4 gnd
port 541 nsew
rlabel metal2 s 15306 3500 15414 3610 4 gnd
port 541 nsew
rlabel metal2 s 2058 14024 2166 14100 4 gnd
port 541 nsew
rlabel metal2 s 15786 25620 15894 25730 4 gnd
port 541 nsew
rlabel metal2 s 18282 11654 18390 11730 4 gnd
port 541 nsew
rlabel metal2 s 810 24610 918 24686 4 gnd
port 541 nsew
rlabel metal2 s 17034 9600 17142 9676 4 gnd
port 541 nsew
rlabel metal2 s 11562 21670 11670 21780 4 gnd
port 541 nsew
rlabel metal2 s 4074 19870 4182 19946 4 gnd
port 541 nsew
rlabel metal2 s 8298 24610 8406 24686 4 gnd
port 541 nsew
rlabel metal2 s 14058 19554 14166 19630 4 gnd
port 541 nsew
rlabel metal2 s 6570 340 6678 450 4 gnd
port 541 nsew
rlabel metal2 s 7050 16930 7158 17040 4 gnd
port 541 nsew
rlabel metal2 s 5802 11654 5910 11730 4 gnd
port 541 nsew
rlabel metal2 s 17034 14024 17142 14100 4 gnd
port 541 nsew
rlabel metal2 s 19050 18290 19158 18366 4 gnd
port 541 nsew
rlabel metal2 s 2058 21450 2166 21526 4 gnd
port 541 nsew
rlabel metal2 s 10314 4544 10422 4620 4 gnd
port 541 nsew
rlabel metal2 s 19050 14340 19158 14416 4 gnd
port 541 nsew
rlabel metal2 s 810 9600 918 9676 4 gnd
port 541 nsew
rlabel metal2 s 18282 9030 18390 9140 4 gnd
port 541 nsew
rlabel metal2 s 12810 16710 12918 16786 4 gnd
port 541 nsew
rlabel metal2 s 9546 17500 9654 17576 4 gnd
port 541 nsew
rlabel metal2 s 13290 10610 13398 10720 4 gnd
port 541 nsew
rlabel metal2 s 20778 340 20886 450 4 gnd
port 541 nsew
rlabel metal2 s 19530 5080 19638 5190 4 gnd
port 541 nsew
rlabel metal2 s 12810 11400 12918 11510 4 gnd
port 541 nsew
rlabel metal2 s 810 13770 918 13880 4 gnd
port 541 nsew
rlabel metal2 s 15786 24294 15894 24370 4 gnd
port 541 nsew
rlabel metal2 s 15786 8810 15894 8886 4 gnd
port 541 nsew
rlabel metal2 s 3306 11654 3414 11730 4 gnd
port 541 nsew
rlabel metal2 s 17802 3754 17910 3830 4 gnd
port 541 nsew
rlabel metal2 s 15786 12444 15894 12520 4 gnd
port 541 nsew
rlabel metal2 s 5802 14024 5910 14100 4 gnd
port 541 nsew
rlabel metal2 s 2826 2490 2934 2566 4 gnd
port 541 nsew
rlabel metal2 s 4554 11400 4662 11510 4 gnd
port 541 nsew
rlabel metal2 s 2826 8020 2934 8096 4 gnd
port 541 nsew
rlabel metal2 s 9066 120 9174 196 4 gnd
port 541 nsew
rlabel metal2 s 6570 22460 6678 22570 4 gnd
port 541 nsew
rlabel metal2 s 10794 594 10902 670 4 gnd
port 541 nsew
rlabel metal2 s 11562 8494 11670 8570 4 gnd
port 541 nsew
rlabel metal2 s 330 12190 438 12300 4 gnd
port 541 nsew
rlabel metal2 s 17034 19870 17142 19946 4 gnd
port 541 nsew
rlabel metal2 s 20778 12444 20886 12520 4 gnd
port 541 nsew
rlabel metal2 s 10314 21670 10422 21780 4 gnd
port 541 nsew
rlabel metal2 s 14538 23820 14646 23896 4 gnd
port 541 nsew
rlabel metal2 s 5802 25084 5910 25160 4 gnd
port 541 nsew
rlabel metal2 s 15786 5080 15894 5190 4 gnd
port 541 nsew
rlabel metal2 s 20778 910 20886 986 4 gnd
port 541 nsew
rlabel metal2 s 12042 18764 12150 18840 4 gnd
port 541 nsew
rlabel metal2 s 10314 8020 10422 8096 4 gnd
port 541 nsew
rlabel metal2 s 14058 7704 14166 7780 4 gnd
port 541 nsew
rlabel metal2 s 11562 16710 11670 16786 4 gnd
port 541 nsew
rlabel metal2 s 9066 6124 9174 6200 4 gnd
port 541 nsew
rlabel metal2 s 19530 9820 19638 9930 4 gnd
port 541 nsew
rlabel metal2 s 7050 11654 7158 11730 4 gnd
port 541 nsew
rlabel metal2 s 19050 3280 19158 3356 4 gnd
port 541 nsew
rlabel metal2 s 19050 19870 19158 19946 4 gnd
port 541 nsew
rlabel metal2 s 16554 2964 16662 3040 4 gnd
port 541 nsew
rlabel metal2 s 4554 3280 4662 3356 4 gnd
port 541 nsew
rlabel metal2 s 3306 21134 3414 21210 4 gnd
port 541 nsew
rlabel metal2 s 16554 3754 16662 3830 4 gnd
port 541 nsew
rlabel metal2 s 12042 23504 12150 23580 4 gnd
port 541 nsew
rlabel metal2 s 12810 11970 12918 12046 4 gnd
port 541 nsew
rlabel metal2 s 12042 3280 12150 3356 4 gnd
port 541 nsew
rlabel metal2 s 17802 25400 17910 25476 4 gnd
port 541 nsew
rlabel metal2 s 12042 7450 12150 7560 4 gnd
port 541 nsew
rlabel metal2 s 13290 6660 13398 6770 4 gnd
port 541 nsew
rlabel metal2 s 3306 6440 3414 6516 4 gnd
port 541 nsew
rlabel metal2 s 7050 8494 7158 8570 4 gnd
port 541 nsew
rlabel metal2 s 12810 17720 12918 17830 4 gnd
port 541 nsew
rlabel metal2 s 9546 10074 9654 10150 4 gnd
port 541 nsew
rlabel metal2 s 20778 6914 20886 6990 4 gnd
port 541 nsew
rlabel metal2 s 5322 9600 5430 9676 4 gnd
port 541 nsew
rlabel metal2 s 4074 4544 4182 4620 4 gnd
port 541 nsew
rlabel metal2 s 15306 1130 15414 1240 4 gnd
port 541 nsew
rlabel metal2 s 9546 15604 9654 15680 4 gnd
port 541 nsew
rlabel metal2 s 330 24040 438 24150 4 gnd
port 541 nsew
rlabel metal2 s 19050 15920 19158 15996 4 gnd
port 541 nsew
rlabel metal2 s 14538 11970 14646 12046 4 gnd
port 541 nsew
rlabel metal2 s 330 23820 438 23896 4 gnd
port 541 nsew
rlabel metal2 s 6570 19080 6678 19156 4 gnd
port 541 nsew
rlabel metal2 s 11562 16930 11670 17040 4 gnd
port 541 nsew
rlabel metal2 s 10794 24040 10902 24150 4 gnd
port 541 nsew
rlabel metal2 s 11562 5334 11670 5410 4 gnd
port 541 nsew
rlabel metal2 s 15786 6660 15894 6770 4 gnd
port 541 nsew
rlabel metal2 s 5322 13550 5430 13626 4 gnd
port 541 nsew
rlabel metal2 s 17802 9600 17910 9676 4 gnd
port 541 nsew
rlabel metal2 s 2058 1130 2166 1240 4 gnd
port 541 nsew
rlabel metal2 s 19530 21924 19638 22000 4 gnd
port 541 nsew
rlabel metal2 s 19530 2964 19638 3040 4 gnd
port 541 nsew
rlabel metal2 s 13290 7704 13398 7780 4 gnd
port 541 nsew
rlabel metal2 s 9546 6660 9654 6770 4 gnd
port 541 nsew
rlabel metal2 s 7050 14814 7158 14890 4 gnd
port 541 nsew
rlabel metal2 s 4074 12760 4182 12836 4 gnd
port 541 nsew
rlabel metal2 s 2826 8494 2934 8570 4 gnd
port 541 nsew
rlabel metal2 s 10794 6440 10902 6516 4 gnd
port 541 nsew
rlabel metal2 s 15786 6440 15894 6516 4 gnd
port 541 nsew
rlabel metal2 s 12810 5650 12918 5726 4 gnd
port 541 nsew
rlabel metal2 s 810 12980 918 13090 4 gnd
port 541 nsew
rlabel metal2 s 14538 19870 14646 19946 4 gnd
port 541 nsew
rlabel metal2 s 20298 18290 20406 18366 4 gnd
port 541 nsew
rlabel metal2 s 19530 14560 19638 14670 4 gnd
port 541 nsew
rlabel metal2 s 9546 15350 9654 15460 4 gnd
port 541 nsew
rlabel metal2 s 10314 340 10422 450 4 gnd
port 541 nsew
rlabel metal2 s 12810 11654 12918 11730 4 gnd
port 541 nsew
rlabel metal2 s 5322 19870 5430 19946 4 gnd
port 541 nsew
rlabel metal2 s 330 8494 438 8570 4 gnd
port 541 nsew
rlabel metal2 s 16554 7450 16662 7560 4 gnd
port 541 nsew
rlabel metal2 s 9546 12190 9654 12300 4 gnd
port 541 nsew
rlabel metal2 s 1578 19300 1686 19410 4 gnd
port 541 nsew
rlabel metal2 s 9066 6914 9174 6990 4 gnd
port 541 nsew
rlabel metal2 s 16554 24040 16662 24150 4 gnd
port 541 nsew
rlabel metal2 s 12810 19554 12918 19630 4 gnd
port 541 nsew
rlabel metal2 s 14538 12980 14646 13090 4 gnd
port 541 nsew
rlabel metal2 s 18282 16140 18390 16250 4 gnd
port 541 nsew
rlabel metal2 s 9066 11180 9174 11256 4 gnd
port 541 nsew
rlabel metal2 s 5322 18510 5430 18620 4 gnd
port 541 nsew
rlabel metal2 s 17034 7704 17142 7780 4 gnd
port 541 nsew
rlabel metal2 s 19530 12444 19638 12520 4 gnd
port 541 nsew
rlabel metal2 s 18282 14814 18390 14890 4 gnd
port 541 nsew
rlabel metal2 s 20298 1384 20406 1460 4 gnd
port 541 nsew
rlabel metal2 s 4554 22460 4662 22570 4 gnd
port 541 nsew
rlabel metal2 s 19530 7230 19638 7306 4 gnd
port 541 nsew
rlabel metal2 s 10314 9820 10422 9930 4 gnd
port 541 nsew
rlabel metal2 s 330 15350 438 15460 4 gnd
port 541 nsew
rlabel metal2 s 4074 9820 4182 9930 4 gnd
port 541 nsew
rlabel metal2 s 5322 14024 5430 14100 4 gnd
port 541 nsew
rlabel metal2 s 9066 3754 9174 3830 4 gnd
port 541 nsew
rlabel metal2 s 8298 23820 8406 23896 4 gnd
port 541 nsew
rlabel metal2 s 19050 9600 19158 9676 4 gnd
port 541 nsew
rlabel metal2 s 5802 910 5910 986 4 gnd
port 541 nsew
rlabel metal2 s 14058 14024 14166 14100 4 gnd
port 541 nsew
rlabel metal2 s 7818 13234 7926 13310 4 gnd
port 541 nsew
rlabel metal2 s 17034 24040 17142 24150 4 gnd
port 541 nsew
rlabel metal2 s 12810 15604 12918 15680 4 gnd
port 541 nsew
rlabel metal2 s 17802 19870 17910 19946 4 gnd
port 541 nsew
rlabel metal2 s 9546 22460 9654 22570 4 gnd
port 541 nsew
rlabel metal2 s 2058 20344 2166 20420 4 gnd
port 541 nsew
rlabel metal2 s 20298 9030 20406 9140 4 gnd
port 541 nsew
rlabel metal2 s 20298 7230 20406 7306 4 gnd
port 541 nsew
rlabel metal2 s 330 2964 438 3040 4 gnd
port 541 nsew
rlabel metal2 s 12042 24830 12150 24940 4 gnd
port 541 nsew
rlabel metal2 s 9066 24294 9174 24370 4 gnd
port 541 nsew
rlabel metal2 s 10794 15130 10902 15206 4 gnd
port 541 nsew
rlabel metal2 s 20778 13550 20886 13626 4 gnd
port 541 nsew
rlabel metal2 s 9066 13234 9174 13310 4 gnd
port 541 nsew
rlabel metal2 s 6570 4070 6678 4146 4 gnd
port 541 nsew
rlabel metal2 s 7818 9030 7926 9140 4 gnd
port 541 nsew
rlabel metal2 s 7818 5650 7926 5726 4 gnd
port 541 nsew
rlabel metal2 s 1578 8240 1686 8350 4 gnd
port 541 nsew
rlabel metal2 s 10794 12444 10902 12520 4 gnd
port 541 nsew
rlabel metal2 s 14058 11654 14166 11730 4 gnd
port 541 nsew
rlabel metal2 s 17802 15130 17910 15206 4 gnd
port 541 nsew
rlabel metal2 s 4074 15920 4182 15996 4 gnd
port 541 nsew
rlabel metal2 s 1578 340 1686 450 4 gnd
port 541 nsew
rlabel metal2 s 4074 1920 4182 2030 4 gnd
port 541 nsew
rlabel metal2 s 17802 23030 17910 23106 4 gnd
port 541 nsew
rlabel metal2 s 7818 16140 7926 16250 4 gnd
port 541 nsew
rlabel metal2 s 330 4860 438 4936 4 gnd
port 541 nsew
rlabel metal2 s 8298 13550 8406 13626 4 gnd
port 541 nsew
rlabel metal2 s 18282 25620 18390 25730 4 gnd
port 541 nsew
rlabel metal2 s 14058 340 14166 450 4 gnd
port 541 nsew
rlabel metal2 s 12810 9030 12918 9140 4 gnd
port 541 nsew
rlabel metal2 s 16554 2490 16662 2566 4 gnd
port 541 nsew
rlabel metal2 s 14058 9284 14166 9360 4 gnd
port 541 nsew
rlabel metal2 s 7818 1384 7926 1460 4 gnd
port 541 nsew
rlabel metal2 s 14538 25400 14646 25476 4 gnd
port 541 nsew
rlabel metal2 s 7050 22240 7158 22316 4 gnd
port 541 nsew
rlabel metal2 s 2058 20880 2166 20990 4 gnd
port 541 nsew
rlabel metal2 s 16554 5334 16662 5410 4 gnd
port 541 nsew
rlabel metal2 s 11562 15920 11670 15996 4 gnd
port 541 nsew
rlabel metal2 s 6570 20344 6678 20420 4 gnd
port 541 nsew
rlabel metal2 s 5322 12980 5430 13090 4 gnd
port 541 nsew
rlabel metal2 s 330 4290 438 4400 4 gnd
port 541 nsew
rlabel metal2 s 2058 23250 2166 23360 4 gnd
port 541 nsew
rlabel metal2 s 18282 12760 18390 12836 4 gnd
port 541 nsew
rlabel metal2 s 12042 7230 12150 7306 4 gnd
port 541 nsew
rlabel metal2 s 7818 19300 7926 19410 4 gnd
port 541 nsew
rlabel metal2 s 3306 13234 3414 13310 4 gnd
port 541 nsew
rlabel metal2 s 17034 10074 17142 10150 4 gnd
port 541 nsew
rlabel metal2 s 7050 3500 7158 3610 4 gnd
port 541 nsew
rlabel metal2 s 5322 9030 5430 9140 4 gnd
port 541 nsew
rlabel metal2 s 20298 1130 20406 1240 4 gnd
port 541 nsew
rlabel metal2 s 19050 12980 19158 13090 4 gnd
port 541 nsew
rlabel metal2 s 5322 13770 5430 13880 4 gnd
port 541 nsew
rlabel metal2 s 2826 16930 2934 17040 4 gnd
port 541 nsew
rlabel metal2 s 4074 25874 4182 25950 4 gnd
port 541 nsew
rlabel metal2 s 9546 21134 9654 21210 4 gnd
port 541 nsew
rlabel metal2 s 20778 13234 20886 13310 4 gnd
port 541 nsew
rlabel metal2 s 11562 21450 11670 21526 4 gnd
port 541 nsew
rlabel metal2 s 20778 17720 20886 17830 4 gnd
port 541 nsew
rlabel metal2 s 5322 10390 5430 10466 4 gnd
port 541 nsew
rlabel metal2 s 12810 2490 12918 2566 4 gnd
port 541 nsew
rlabel metal2 s 20298 10390 20406 10466 4 gnd
port 541 nsew
rlabel metal2 s 2826 8810 2934 8886 4 gnd
port 541 nsew
rlabel metal2 s 2826 7704 2934 7780 4 gnd
port 541 nsew
rlabel metal2 s 9546 11180 9654 11256 4 gnd
port 541 nsew
rlabel metal2 s 2058 5870 2166 5980 4 gnd
port 541 nsew
rlabel metal2 s 18282 9820 18390 9930 4 gnd
port 541 nsew
rlabel metal2 s 15786 2174 15894 2250 4 gnd
port 541 nsew
rlabel metal2 s 7818 14814 7926 14890 4 gnd
port 541 nsew
rlabel metal2 s 20298 9284 20406 9360 4 gnd
port 541 nsew
rlabel metal2 s 17802 120 17910 196 4 gnd
port 541 nsew
rlabel metal2 s 17034 9030 17142 9140 4 gnd
port 541 nsew
rlabel metal2 s 4554 2710 4662 2820 4 gnd
port 541 nsew
rlabel metal2 s 13290 20880 13398 20990 4 gnd
port 541 nsew
rlabel metal2 s 15786 3280 15894 3356 4 gnd
port 541 nsew
rlabel metal2 s 15786 21924 15894 22000 4 gnd
port 541 nsew
rlabel metal2 s 10314 12444 10422 12520 4 gnd
port 541 nsew
rlabel metal2 s 19530 1700 19638 1776 4 gnd
port 541 nsew
rlabel metal2 s 17802 23504 17910 23580 4 gnd
port 541 nsew
rlabel metal2 s 10314 24040 10422 24150 4 gnd
port 541 nsew
rlabel metal2 s 11562 21134 11670 21210 4 gnd
port 541 nsew
rlabel metal2 s 4554 9284 4662 9360 4 gnd
port 541 nsew
rlabel metal2 s 15786 120 15894 196 4 gnd
port 541 nsew
rlabel metal2 s 16554 16394 16662 16470 4 gnd
port 541 nsew
rlabel metal2 s 14058 9600 14166 9676 4 gnd
port 541 nsew
rlabel metal2 s 10794 6124 10902 6200 4 gnd
port 541 nsew
rlabel metal2 s 20778 24610 20886 24686 4 gnd
port 541 nsew
rlabel metal2 s 18282 21924 18390 22000 4 gnd
port 541 nsew
rlabel metal2 s 9066 17720 9174 17830 4 gnd
port 541 nsew
rlabel metal2 s 17802 13770 17910 13880 4 gnd
port 541 nsew
rlabel metal2 s 6570 21670 6678 21780 4 gnd
port 541 nsew
rlabel metal2 s 13290 18290 13398 18366 4 gnd
port 541 nsew
rlabel metal2 s 12042 4544 12150 4620 4 gnd
port 541 nsew
rlabel metal2 s 330 19554 438 19630 4 gnd
port 541 nsew
rlabel metal2 s 330 9030 438 9140 4 gnd
port 541 nsew
rlabel metal2 s 12042 25400 12150 25476 4 gnd
port 541 nsew
rlabel metal2 s 10794 3500 10902 3610 4 gnd
port 541 nsew
rlabel metal2 s 20298 17500 20406 17576 4 gnd
port 541 nsew
rlabel metal2 s 6570 8240 6678 8350 4 gnd
port 541 nsew
rlabel metal2 s 16554 21670 16662 21780 4 gnd
port 541 nsew
rlabel metal2 s 14058 21134 14166 21210 4 gnd
port 541 nsew
rlabel metal2 s 13290 21670 13398 21780 4 gnd
port 541 nsew
rlabel metal2 s 19050 12760 19158 12836 4 gnd
port 541 nsew
rlabel metal2 s 12042 1130 12150 1240 4 gnd
port 541 nsew
rlabel metal2 s 19050 8494 19158 8570 4 gnd
port 541 nsew
rlabel metal2 s 4074 19080 4182 19156 4 gnd
port 541 nsew
rlabel metal2 s 6570 21924 6678 22000 4 gnd
port 541 nsew
rlabel metal2 s 12810 21450 12918 21526 4 gnd
port 541 nsew
rlabel metal2 s 8298 25620 8406 25730 4 gnd
port 541 nsew
rlabel metal2 s 8298 15130 8406 15206 4 gnd
port 541 nsew
rlabel metal2 s 15786 25084 15894 25160 4 gnd
port 541 nsew
rlabel metal2 s 9546 23504 9654 23580 4 gnd
port 541 nsew
rlabel metal2 s 5322 24294 5430 24370 4 gnd
port 541 nsew
rlabel metal2 s 7050 22714 7158 22790 4 gnd
port 541 nsew
rlabel metal2 s 20778 5334 20886 5410 4 gnd
port 541 nsew
rlabel metal2 s 9066 12190 9174 12300 4 gnd
port 541 nsew
rlabel metal2 s 1578 23820 1686 23896 4 gnd
port 541 nsew
rlabel metal2 s 20778 2710 20886 2820 4 gnd
port 541 nsew
rlabel metal2 s 11562 16140 11670 16250 4 gnd
port 541 nsew
rlabel metal2 s 17802 10864 17910 10940 4 gnd
port 541 nsew
rlabel metal2 s 13290 13234 13398 13310 4 gnd
port 541 nsew
rlabel metal2 s 20298 19554 20406 19630 4 gnd
port 541 nsew
rlabel metal2 s 810 22714 918 22790 4 gnd
port 541 nsew
rlabel metal2 s 4074 8494 4182 8570 4 gnd
port 541 nsew
rlabel metal2 s 810 3280 918 3356 4 gnd
port 541 nsew
rlabel metal2 s 19530 23250 19638 23360 4 gnd
port 541 nsew
rlabel metal2 s 15786 25874 15894 25950 4 gnd
port 541 nsew
rlabel metal2 s 15306 8810 15414 8886 4 gnd
port 541 nsew
rlabel metal2 s 11562 4070 11670 4146 4 gnd
port 541 nsew
rlabel metal2 s 15786 17974 15894 18050 4 gnd
port 541 nsew
rlabel metal2 s 810 1920 918 2030 4 gnd
port 541 nsew
rlabel metal2 s 11562 21924 11670 22000 4 gnd
port 541 nsew
rlabel metal2 s 11562 23030 11670 23106 4 gnd
port 541 nsew
rlabel metal2 s 5322 22460 5430 22570 4 gnd
port 541 nsew
rlabel metal2 s 8298 25400 8406 25476 4 gnd
port 541 nsew
rlabel metal2 s 18282 25400 18390 25476 4 gnd
port 541 nsew
rlabel metal2 s 8298 14560 8406 14670 4 gnd
port 541 nsew
rlabel metal2 s 12810 25874 12918 25950 4 gnd
port 541 nsew
rlabel metal2 s 14538 1700 14646 1776 4 gnd
port 541 nsew
rlabel metal2 s 18282 8494 18390 8570 4 gnd
port 541 nsew
rlabel metal2 s 810 10610 918 10720 4 gnd
port 541 nsew
rlabel metal2 s 9066 5650 9174 5726 4 gnd
port 541 nsew
rlabel metal2 s 18282 15920 18390 15996 4 gnd
port 541 nsew
rlabel metal2 s 17802 21924 17910 22000 4 gnd
port 541 nsew
rlabel metal2 s 19050 21134 19158 21210 4 gnd
port 541 nsew
rlabel metal2 s 1578 5650 1686 5726 4 gnd
port 541 nsew
rlabel metal2 s 16554 19080 16662 19156 4 gnd
port 541 nsew
rlabel metal2 s 9546 24294 9654 24370 4 gnd
port 541 nsew
rlabel metal2 s 6570 7704 6678 7780 4 gnd
port 541 nsew
rlabel metal2 s 4554 10390 4662 10466 4 gnd
port 541 nsew
rlabel metal2 s 3306 20344 3414 20420 4 gnd
port 541 nsew
rlabel metal2 s 9546 9284 9654 9360 4 gnd
port 541 nsew
rlabel metal2 s 9546 1384 9654 1460 4 gnd
port 541 nsew
rlabel metal2 s 810 20660 918 20736 4 gnd
port 541 nsew
rlabel metal2 s 2058 18510 2166 18620 4 gnd
port 541 nsew
rlabel metal2 s 10794 12760 10902 12836 4 gnd
port 541 nsew
rlabel metal2 s 14058 17184 14166 17260 4 gnd
port 541 nsew
rlabel metal2 s 7050 18290 7158 18366 4 gnd
port 541 nsew
rlabel metal2 s 810 3754 918 3830 4 gnd
port 541 nsew
rlabel metal2 s 16554 10864 16662 10940 4 gnd
port 541 nsew
rlabel metal2 s 6570 6914 6678 6990 4 gnd
port 541 nsew
rlabel metal2 s 20778 23820 20886 23896 4 gnd
port 541 nsew
rlabel metal2 s 19530 22240 19638 22316 4 gnd
port 541 nsew
rlabel metal2 s 18282 10074 18390 10150 4 gnd
port 541 nsew
rlabel metal2 s 2058 8810 2166 8886 4 gnd
port 541 nsew
rlabel metal2 s 7818 25084 7926 25160 4 gnd
port 541 nsew
rlabel metal2 s 11562 1384 11670 1460 4 gnd
port 541 nsew
rlabel metal2 s 7050 19080 7158 19156 4 gnd
port 541 nsew
rlabel metal2 s 810 15920 918 15996 4 gnd
port 541 nsew
rlabel metal2 s 7050 6124 7158 6200 4 gnd
port 541 nsew
rlabel metal2 s 1578 3280 1686 3356 4 gnd
port 541 nsew
rlabel metal2 s 17034 21924 17142 22000 4 gnd
port 541 nsew
rlabel metal2 s 2826 14340 2934 14416 4 gnd
port 541 nsew
rlabel metal2 s 5322 25400 5430 25476 4 gnd
port 541 nsew
rlabel metal2 s 330 18290 438 18366 4 gnd
port 541 nsew
rlabel metal2 s 10794 5334 10902 5410 4 gnd
port 541 nsew
rlabel metal2 s 8298 2964 8406 3040 4 gnd
port 541 nsew
rlabel metal2 s 20778 16140 20886 16250 4 gnd
port 541 nsew
rlabel metal2 s 810 8810 918 8886 4 gnd
port 541 nsew
rlabel metal2 s 6570 23504 6678 23580 4 gnd
port 541 nsew
rlabel metal2 s 810 6660 918 6770 4 gnd
port 541 nsew
rlabel metal2 s 810 16140 918 16250 4 gnd
port 541 nsew
rlabel metal2 s 12042 20660 12150 20736 4 gnd
port 541 nsew
rlabel metal2 s 12810 1130 12918 1240 4 gnd
port 541 nsew
rlabel metal2 s 11562 10610 11670 10720 4 gnd
port 541 nsew
rlabel metal2 s 14058 1384 14166 1460 4 gnd
port 541 nsew
rlabel metal2 s 12810 7230 12918 7306 4 gnd
port 541 nsew
rlabel metal2 s 17802 25874 17910 25950 4 gnd
port 541 nsew
rlabel metal2 s 4074 16930 4182 17040 4 gnd
port 541 nsew
rlabel metal2 s 10794 8494 10902 8570 4 gnd
port 541 nsew
rlabel metal2 s 20778 2964 20886 3040 4 gnd
port 541 nsew
rlabel metal2 s 10794 9600 10902 9676 4 gnd
port 541 nsew
rlabel metal2 s 1578 7704 1686 7780 4 gnd
port 541 nsew
rlabel metal2 s 15786 14024 15894 14100 4 gnd
port 541 nsew
rlabel metal2 s 19050 9820 19158 9930 4 gnd
port 541 nsew
rlabel metal2 s 13290 2490 13398 2566 4 gnd
port 541 nsew
rlabel metal2 s 10314 8240 10422 8350 4 gnd
port 541 nsew
rlabel metal2 s 7818 23820 7926 23896 4 gnd
port 541 nsew
rlabel metal2 s 810 6124 918 6200 4 gnd
port 541 nsew
rlabel metal2 s 17034 17720 17142 17830 4 gnd
port 541 nsew
rlabel metal2 s 17034 20090 17142 20200 4 gnd
port 541 nsew
rlabel metal2 s 7818 8810 7926 8886 4 gnd
port 541 nsew
rlabel metal2 s 6570 19300 6678 19410 4 gnd
port 541 nsew
rlabel metal2 s 4554 120 4662 196 4 gnd
port 541 nsew
rlabel metal2 s 9546 12444 9654 12520 4 gnd
port 541 nsew
rlabel metal2 s 3306 9030 3414 9140 4 gnd
port 541 nsew
rlabel metal2 s 5322 9284 5430 9360 4 gnd
port 541 nsew
rlabel metal2 s 13290 15350 13398 15460 4 gnd
port 541 nsew
rlabel metal2 s 2058 16710 2166 16786 4 gnd
port 541 nsew
rlabel metal2 s 17034 21670 17142 21780 4 gnd
port 541 nsew
rlabel metal2 s 12042 16394 12150 16470 4 gnd
port 541 nsew
rlabel metal2 s 4554 14814 4662 14890 4 gnd
port 541 nsew
rlabel metal2 s 2826 19080 2934 19156 4 gnd
port 541 nsew
rlabel metal2 s 5802 12760 5910 12836 4 gnd
port 541 nsew
rlabel metal2 s 18282 1700 18390 1776 4 gnd
port 541 nsew
rlabel metal2 s 17034 8240 17142 8350 4 gnd
port 541 nsew
rlabel metal2 s 9066 340 9174 450 4 gnd
port 541 nsew
rlabel metal2 s 12042 24040 12150 24150 4 gnd
port 541 nsew
rlabel metal2 s 9066 25400 9174 25476 4 gnd
port 541 nsew
rlabel metal2 s 17802 24040 17910 24150 4 gnd
port 541 nsew
rlabel metal2 s 11562 24830 11670 24940 4 gnd
port 541 nsew
rlabel metal2 s 17802 18290 17910 18366 4 gnd
port 541 nsew
rlabel metal2 s 10314 6660 10422 6770 4 gnd
port 541 nsew
rlabel metal2 s 2058 13234 2166 13310 4 gnd
port 541 nsew
rlabel metal2 s 5802 15604 5910 15680 4 gnd
port 541 nsew
rlabel metal2 s 17802 14814 17910 14890 4 gnd
port 541 nsew
rlabel metal2 s 8298 7704 8406 7780 4 gnd
port 541 nsew
rlabel metal2 s 6570 3280 6678 3356 4 gnd
port 541 nsew
rlabel metal2 s 10314 19554 10422 19630 4 gnd
port 541 nsew
rlabel metal2 s 14538 1920 14646 2030 4 gnd
port 541 nsew
rlabel metal2 s 7818 23504 7926 23580 4 gnd
port 541 nsew
rlabel metal2 s 10314 13770 10422 13880 4 gnd
port 541 nsew
rlabel metal2 s 12042 21670 12150 21780 4 gnd
port 541 nsew
rlabel metal2 s 7818 6124 7926 6200 4 gnd
port 541 nsew
rlabel metal2 s 13290 9820 13398 9930 4 gnd
port 541 nsew
rlabel metal2 s 5322 19080 5430 19156 4 gnd
port 541 nsew
rlabel metal2 s 10794 7450 10902 7560 4 gnd
port 541 nsew
rlabel metal2 s 5322 17184 5430 17260 4 gnd
port 541 nsew
rlabel metal2 s 7818 24610 7926 24686 4 gnd
port 541 nsew
rlabel metal2 s 5322 910 5430 986 4 gnd
port 541 nsew
rlabel metal2 s 5322 3754 5430 3830 4 gnd
port 541 nsew
rlabel metal2 s 20778 25084 20886 25160 4 gnd
port 541 nsew
rlabel metal2 s 7050 11400 7158 11510 4 gnd
port 541 nsew
rlabel metal2 s 10314 15920 10422 15996 4 gnd
port 541 nsew
rlabel metal2 s 15306 17720 15414 17830 4 gnd
port 541 nsew
rlabel metal2 s 1578 4544 1686 4620 4 gnd
port 541 nsew
rlabel metal2 s 14538 15920 14646 15996 4 gnd
port 541 nsew
rlabel metal2 s 2826 25400 2934 25476 4 gnd
port 541 nsew
rlabel metal2 s 6570 13770 6678 13880 4 gnd
port 541 nsew
rlabel metal2 s 17034 6124 17142 6200 4 gnd
port 541 nsew
rlabel metal2 s 15306 19870 15414 19946 4 gnd
port 541 nsew
rlabel metal2 s 16554 23504 16662 23580 4 gnd
port 541 nsew
rlabel metal2 s 330 12760 438 12836 4 gnd
port 541 nsew
rlabel metal2 s 1578 12760 1686 12836 4 gnd
port 541 nsew
rlabel metal2 s 11562 18764 11670 18840 4 gnd
port 541 nsew
rlabel metal2 s 4074 8020 4182 8096 4 gnd
port 541 nsew
rlabel metal2 s 15786 5334 15894 5410 4 gnd
port 541 nsew
rlabel metal2 s 19530 10074 19638 10150 4 gnd
port 541 nsew
rlabel metal2 s 810 21670 918 21780 4 gnd
port 541 nsew
rlabel metal2 s 4554 9030 4662 9140 4 gnd
port 541 nsew
rlabel metal2 s 5802 19554 5910 19630 4 gnd
port 541 nsew
rlabel metal2 s 6570 22240 6678 22316 4 gnd
port 541 nsew
rlabel metal2 s 10794 21670 10902 21780 4 gnd
port 541 nsew
rlabel metal2 s 19050 6440 19158 6516 4 gnd
port 541 nsew
rlabel metal2 s 1578 25874 1686 25950 4 gnd
port 541 nsew
rlabel metal2 s 19050 24610 19158 24686 4 gnd
port 541 nsew
rlabel metal2 s 10314 8494 10422 8570 4 gnd
port 541 nsew
rlabel metal2 s 7050 19300 7158 19410 4 gnd
port 541 nsew
rlabel metal2 s 10314 21924 10422 22000 4 gnd
port 541 nsew
rlabel metal2 s 3306 5870 3414 5980 4 gnd
port 541 nsew
rlabel metal2 s 9546 20880 9654 20990 4 gnd
port 541 nsew
rlabel metal2 s 10794 16930 10902 17040 4 gnd
port 541 nsew
rlabel metal2 s 10314 7450 10422 7560 4 gnd
port 541 nsew
rlabel metal2 s 15786 18510 15894 18620 4 gnd
port 541 nsew
rlabel metal2 s 15786 5650 15894 5726 4 gnd
port 541 nsew
rlabel metal2 s 16554 6440 16662 6516 4 gnd
port 541 nsew
rlabel metal2 s 18282 6660 18390 6770 4 gnd
port 541 nsew
rlabel metal2 s 9066 23820 9174 23896 4 gnd
port 541 nsew
rlabel metal2 s 6570 4860 6678 4936 4 gnd
port 541 nsew
rlabel metal2 s 19050 1700 19158 1776 4 gnd
port 541 nsew
rlabel metal2 s 19530 8240 19638 8350 4 gnd
port 541 nsew
rlabel metal2 s 17802 20344 17910 20420 4 gnd
port 541 nsew
rlabel metal2 s 17034 16140 17142 16250 4 gnd
port 541 nsew
rlabel metal2 s 7050 1384 7158 1460 4 gnd
port 541 nsew
rlabel metal2 s 17802 7230 17910 7306 4 gnd
port 541 nsew
rlabel metal2 s 15306 9030 15414 9140 4 gnd
port 541 nsew
rlabel metal2 s 5322 15604 5430 15680 4 gnd
port 541 nsew
rlabel metal2 s 16554 22460 16662 22570 4 gnd
port 541 nsew
rlabel metal2 s 6570 16394 6678 16470 4 gnd
port 541 nsew
rlabel metal2 s 2826 12760 2934 12836 4 gnd
port 541 nsew
rlabel metal2 s 9066 8494 9174 8570 4 gnd
port 541 nsew
rlabel metal2 s 14538 11180 14646 11256 4 gnd
port 541 nsew
rlabel metal2 s 3306 9820 3414 9930 4 gnd
port 541 nsew
rlabel metal2 s 17034 23250 17142 23360 4 gnd
port 541 nsew
rlabel metal2 s 19050 15604 19158 15680 4 gnd
port 541 nsew
rlabel metal2 s 15786 18764 15894 18840 4 gnd
port 541 nsew
rlabel metal2 s 5802 6914 5910 6990 4 gnd
port 541 nsew
rlabel metal2 s 15306 2174 15414 2250 4 gnd
port 541 nsew
rlabel metal2 s 810 18764 918 18840 4 gnd
port 541 nsew
rlabel metal2 s 5802 8020 5910 8096 4 gnd
port 541 nsew
rlabel metal2 s 2826 11400 2934 11510 4 gnd
port 541 nsew
rlabel metal2 s 17034 15350 17142 15460 4 gnd
port 541 nsew
rlabel metal2 s 9546 5870 9654 5980 4 gnd
port 541 nsew
rlabel metal2 s 12042 17184 12150 17260 4 gnd
port 541 nsew
rlabel metal2 s 17802 17720 17910 17830 4 gnd
port 541 nsew
rlabel metal2 s 8298 2710 8406 2820 4 gnd
port 541 nsew
rlabel metal2 s 3306 24294 3414 24370 4 gnd
port 541 nsew
rlabel metal2 s 17802 22240 17910 22316 4 gnd
port 541 nsew
rlabel metal2 s 4554 2490 4662 2566 4 gnd
port 541 nsew
rlabel metal2 s 10314 10610 10422 10720 4 gnd
port 541 nsew
rlabel metal2 s 10794 14024 10902 14100 4 gnd
port 541 nsew
rlabel metal2 s 4554 14560 4662 14670 4 gnd
port 541 nsew
rlabel metal2 s 19530 10610 19638 10720 4 gnd
port 541 nsew
rlabel metal2 s 20298 9820 20406 9930 4 gnd
port 541 nsew
rlabel metal2 s 13290 20344 13398 20420 4 gnd
port 541 nsew
rlabel metal2 s 9546 24610 9654 24686 4 gnd
port 541 nsew
rlabel metal2 s 7818 340 7926 450 4 gnd
port 541 nsew
rlabel metal2 s 330 25400 438 25476 4 gnd
port 541 nsew
rlabel metal2 s 6570 3754 6678 3830 4 gnd
port 541 nsew
rlabel metal2 s 19050 24830 19158 24940 4 gnd
port 541 nsew
rlabel metal2 s 4074 14340 4182 14416 4 gnd
port 541 nsew
rlabel metal2 s 20298 3754 20406 3830 4 gnd
port 541 nsew
rlabel metal2 s 9546 25084 9654 25160 4 gnd
port 541 nsew
rlabel metal2 s 14538 4290 14646 4400 4 gnd
port 541 nsew
rlabel metal2 s 15306 18290 15414 18366 4 gnd
port 541 nsew
rlabel metal2 s 10794 13770 10902 13880 4 gnd
port 541 nsew
rlabel metal2 s 7818 12444 7926 12520 4 gnd
port 541 nsew
rlabel metal2 s 7050 16394 7158 16470 4 gnd
port 541 nsew
rlabel metal2 s 2826 6440 2934 6516 4 gnd
port 541 nsew
rlabel metal2 s 2058 9820 2166 9930 4 gnd
port 541 nsew
rlabel metal2 s 14058 11180 14166 11256 4 gnd
port 541 nsew
rlabel metal2 s 7818 10074 7926 10150 4 gnd
port 541 nsew
rlabel metal2 s 9546 6124 9654 6200 4 gnd
port 541 nsew
rlabel metal2 s 7050 5650 7158 5726 4 gnd
port 541 nsew
rlabel metal2 s 5322 11180 5430 11256 4 gnd
port 541 nsew
rlabel metal2 s 12810 15350 12918 15460 4 gnd
port 541 nsew
rlabel metal2 s 17034 11970 17142 12046 4 gnd
port 541 nsew
rlabel metal2 s 19050 13770 19158 13880 4 gnd
port 541 nsew
rlabel metal2 s 11562 25874 11670 25950 4 gnd
port 541 nsew
rlabel metal2 s 7818 15604 7926 15680 4 gnd
port 541 nsew
rlabel metal2 s 12810 4290 12918 4400 4 gnd
port 541 nsew
rlabel metal2 s 18282 13770 18390 13880 4 gnd
port 541 nsew
rlabel metal2 s 16554 594 16662 670 4 gnd
port 541 nsew
rlabel metal2 s 13290 20090 13398 20200 4 gnd
port 541 nsew
rlabel metal2 s 11562 4544 11670 4620 4 gnd
port 541 nsew
rlabel metal2 s 4074 22714 4182 22790 4 gnd
port 541 nsew
rlabel metal2 s 9066 910 9174 986 4 gnd
port 541 nsew
rlabel metal2 s 11562 15350 11670 15460 4 gnd
port 541 nsew
rlabel metal2 s 8298 4544 8406 4620 4 gnd
port 541 nsew
rlabel metal2 s 19530 11400 19638 11510 4 gnd
port 541 nsew
rlabel metal2 s 3306 6660 3414 6770 4 gnd
port 541 nsew
rlabel metal2 s 15786 14814 15894 14890 4 gnd
port 541 nsew
rlabel metal2 s 13290 6124 13398 6200 4 gnd
port 541 nsew
rlabel metal2 s 19530 19554 19638 19630 4 gnd
port 541 nsew
rlabel metal2 s 20298 18510 20406 18620 4 gnd
port 541 nsew
rlabel metal2 s 10314 4070 10422 4146 4 gnd
port 541 nsew
rlabel metal2 s 13290 16394 13398 16470 4 gnd
port 541 nsew
rlabel metal2 s 2826 20660 2934 20736 4 gnd
port 541 nsew
rlabel metal2 s 10794 6660 10902 6770 4 gnd
port 541 nsew
rlabel metal2 s 4554 910 4662 986 4 gnd
port 541 nsew
rlabel metal2 s 19530 11654 19638 11730 4 gnd
port 541 nsew
rlabel metal2 s 20778 2174 20886 2250 4 gnd
port 541 nsew
rlabel metal2 s 1578 11970 1686 12046 4 gnd
port 541 nsew
rlabel metal2 s 9066 3280 9174 3356 4 gnd
port 541 nsew
rlabel metal2 s 1578 3500 1686 3610 4 gnd
port 541 nsew
rlabel metal2 s 5802 3754 5910 3830 4 gnd
port 541 nsew
rlabel metal2 s 5322 25084 5430 25160 4 gnd
port 541 nsew
rlabel metal2 s 17034 22460 17142 22570 4 gnd
port 541 nsew
rlabel metal2 s 20778 15130 20886 15206 4 gnd
port 541 nsew
rlabel metal2 s 11562 11400 11670 11510 4 gnd
port 541 nsew
rlabel metal2 s 18282 17500 18390 17576 4 gnd
port 541 nsew
rlabel metal2 s 4554 12190 4662 12300 4 gnd
port 541 nsew
rlabel metal2 s 10314 2174 10422 2250 4 gnd
port 541 nsew
rlabel metal2 s 17034 5334 17142 5410 4 gnd
port 541 nsew
rlabel metal2 s 9066 21450 9174 21526 4 gnd
port 541 nsew
rlabel metal2 s 15306 20880 15414 20990 4 gnd
port 541 nsew
rlabel metal2 s 16554 5080 16662 5190 4 gnd
port 541 nsew
rlabel metal2 s 10794 18764 10902 18840 4 gnd
port 541 nsew
rlabel metal2 s 2058 5080 2166 5190 4 gnd
port 541 nsew
rlabel metal2 s 16554 6660 16662 6770 4 gnd
port 541 nsew
rlabel metal2 s 4554 15604 4662 15680 4 gnd
port 541 nsew
rlabel metal2 s 2058 16394 2166 16470 4 gnd
port 541 nsew
rlabel metal2 s 12042 19870 12150 19946 4 gnd
port 541 nsew
rlabel metal2 s 5322 17720 5430 17830 4 gnd
port 541 nsew
rlabel metal2 s 18282 4860 18390 4936 4 gnd
port 541 nsew
rlabel metal2 s 2058 1920 2166 2030 4 gnd
port 541 nsew
rlabel metal2 s 14538 20660 14646 20736 4 gnd
port 541 nsew
rlabel metal2 s 8298 10390 8406 10466 4 gnd
port 541 nsew
rlabel metal2 s 330 16140 438 16250 4 gnd
port 541 nsew
rlabel metal2 s 2058 20090 2166 20200 4 gnd
port 541 nsew
rlabel metal2 s 14538 4860 14646 4936 4 gnd
port 541 nsew
rlabel metal2 s 7050 24040 7158 24150 4 gnd
port 541 nsew
rlabel metal2 s 8298 13234 8406 13310 4 gnd
port 541 nsew
rlabel metal2 s 17034 2710 17142 2820 4 gnd
port 541 nsew
rlabel metal2 s 12810 17974 12918 18050 4 gnd
port 541 nsew
rlabel metal2 s 7050 13770 7158 13880 4 gnd
port 541 nsew
rlabel metal2 s 4554 18290 4662 18366 4 gnd
port 541 nsew
rlabel metal2 s 13290 6440 13398 6516 4 gnd
port 541 nsew
rlabel metal2 s 7050 11970 7158 12046 4 gnd
port 541 nsew
rlabel metal2 s 15786 21670 15894 21780 4 gnd
port 541 nsew
rlabel metal2 s 14538 14560 14646 14670 4 gnd
port 541 nsew
rlabel metal2 s 1578 14814 1686 14890 4 gnd
port 541 nsew
rlabel metal2 s 7818 25874 7926 25950 4 gnd
port 541 nsew
rlabel metal2 s 10314 5334 10422 5410 4 gnd
port 541 nsew
rlabel metal2 s 3306 20660 3414 20736 4 gnd
port 541 nsew
rlabel metal2 s 9066 9600 9174 9676 4 gnd
port 541 nsew
rlabel metal2 s 16554 25400 16662 25476 4 gnd
port 541 nsew
rlabel metal2 s 11562 19554 11670 19630 4 gnd
port 541 nsew
rlabel metal2 s 1578 10864 1686 10940 4 gnd
port 541 nsew
rlabel metal2 s 4554 25400 4662 25476 4 gnd
port 541 nsew
rlabel metal2 s 2058 17500 2166 17576 4 gnd
port 541 nsew
rlabel metal2 s 14538 2964 14646 3040 4 gnd
port 541 nsew
rlabel metal2 s 15786 12190 15894 12300 4 gnd
port 541 nsew
rlabel metal2 s 9066 11400 9174 11510 4 gnd
port 541 nsew
rlabel metal2 s 2826 14560 2934 14670 4 gnd
port 541 nsew
rlabel metal2 s 10794 20344 10902 20420 4 gnd
port 541 nsew
rlabel metal2 s 14538 16710 14646 16786 4 gnd
port 541 nsew
rlabel metal2 s 9066 25874 9174 25950 4 gnd
port 541 nsew
rlabel metal2 s 7050 6660 7158 6770 4 gnd
port 541 nsew
rlabel metal2 s 18282 25084 18390 25160 4 gnd
port 541 nsew
rlabel metal2 s 19530 6124 19638 6200 4 gnd
port 541 nsew
rlabel metal2 s 20298 13770 20406 13880 4 gnd
port 541 nsew
rlabel metal2 s 7818 9284 7926 9360 4 gnd
port 541 nsew
rlabel metal2 s 4074 18510 4182 18620 4 gnd
port 541 nsew
rlabel metal2 s 5322 23250 5430 23360 4 gnd
port 541 nsew
rlabel metal2 s 4554 12760 4662 12836 4 gnd
port 541 nsew
rlabel metal2 s 6570 2174 6678 2250 4 gnd
port 541 nsew
rlabel metal2 s 17802 24830 17910 24940 4 gnd
port 541 nsew
rlabel metal2 s 10794 2490 10902 2566 4 gnd
port 541 nsew
rlabel metal2 s 11562 3754 11670 3830 4 gnd
port 541 nsew
rlabel metal2 s 9066 2490 9174 2566 4 gnd
port 541 nsew
rlabel metal2 s 15306 15350 15414 15460 4 gnd
port 541 nsew
rlabel metal2 s 15306 10864 15414 10940 4 gnd
port 541 nsew
rlabel metal2 s 4074 11400 4182 11510 4 gnd
port 541 nsew
rlabel metal2 s 2058 12190 2166 12300 4 gnd
port 541 nsew
rlabel metal2 s 17034 8020 17142 8096 4 gnd
port 541 nsew
rlabel metal2 s 1578 14024 1686 14100 4 gnd
port 541 nsew
rlabel metal2 s 330 20880 438 20990 4 gnd
port 541 nsew
rlabel metal2 s 15786 2964 15894 3040 4 gnd
port 541 nsew
rlabel metal2 s 17802 16394 17910 16470 4 gnd
port 541 nsew
rlabel metal2 s 8298 19300 8406 19410 4 gnd
port 541 nsew
rlabel metal2 s 14538 13550 14646 13626 4 gnd
port 541 nsew
rlabel metal2 s 16554 14024 16662 14100 4 gnd
port 541 nsew
rlabel metal2 s 4074 23030 4182 23106 4 gnd
port 541 nsew
rlabel metal2 s 1578 9284 1686 9360 4 gnd
port 541 nsew
rlabel metal2 s 19530 17720 19638 17830 4 gnd
port 541 nsew
rlabel metal2 s 6570 13550 6678 13626 4 gnd
port 541 nsew
rlabel metal2 s 2826 14024 2934 14100 4 gnd
port 541 nsew
rlabel metal2 s 7818 12980 7926 13090 4 gnd
port 541 nsew
rlabel metal2 s 8298 18290 8406 18366 4 gnd
port 541 nsew
rlabel metal2 s 10794 4544 10902 4620 4 gnd
port 541 nsew
rlabel metal2 s 18282 15130 18390 15206 4 gnd
port 541 nsew
rlabel metal2 s 4554 24830 4662 24940 4 gnd
port 541 nsew
rlabel metal2 s 13290 12444 13398 12520 4 gnd
port 541 nsew
rlabel metal2 s 19530 1920 19638 2030 4 gnd
port 541 nsew
rlabel metal2 s 7818 910 7926 986 4 gnd
port 541 nsew
rlabel metal2 s 810 15350 918 15460 4 gnd
port 541 nsew
rlabel metal2 s 20298 23030 20406 23106 4 gnd
port 541 nsew
rlabel metal2 s 6570 22714 6678 22790 4 gnd
port 541 nsew
rlabel metal2 s 5322 2964 5430 3040 4 gnd
port 541 nsew
rlabel metal2 s 3306 4860 3414 4936 4 gnd
port 541 nsew
rlabel metal2 s 6570 14814 6678 14890 4 gnd
port 541 nsew
rlabel metal2 s 17034 16710 17142 16786 4 gnd
port 541 nsew
rlabel metal2 s 1578 16930 1686 17040 4 gnd
port 541 nsew
rlabel metal2 s 11562 22240 11670 22316 4 gnd
port 541 nsew
rlabel metal2 s 13290 17500 13398 17576 4 gnd
port 541 nsew
rlabel metal2 s 19050 21924 19158 22000 4 gnd
port 541 nsew
rlabel metal2 s 18282 13234 18390 13310 4 gnd
port 541 nsew
rlabel metal2 s 6570 18510 6678 18620 4 gnd
port 541 nsew
rlabel metal2 s 10794 21924 10902 22000 4 gnd
port 541 nsew
rlabel metal2 s 17034 1384 17142 1460 4 gnd
port 541 nsew
rlabel metal2 s 16554 11180 16662 11256 4 gnd
port 541 nsew
rlabel metal2 s 5322 8810 5430 8886 4 gnd
port 541 nsew
rlabel metal2 s 5802 19080 5910 19156 4 gnd
port 541 nsew
rlabel metal2 s 20778 17184 20886 17260 4 gnd
port 541 nsew
rlabel metal2 s 2058 3754 2166 3830 4 gnd
port 541 nsew
rlabel metal2 s 6570 10074 6678 10150 4 gnd
port 541 nsew
rlabel metal2 s 7818 13770 7926 13880 4 gnd
port 541 nsew
rlabel metal2 s 5322 9820 5430 9930 4 gnd
port 541 nsew
rlabel metal2 s 7818 5870 7926 5980 4 gnd
port 541 nsew
rlabel metal2 s 12810 20880 12918 20990 4 gnd
port 541 nsew
rlabel metal2 s 17034 910 17142 986 4 gnd
port 541 nsew
rlabel metal2 s 810 2490 918 2566 4 gnd
port 541 nsew
rlabel metal2 s 5802 25874 5910 25950 4 gnd
port 541 nsew
rlabel metal2 s 7050 6440 7158 6516 4 gnd
port 541 nsew
rlabel metal2 s 7818 3500 7926 3610 4 gnd
port 541 nsew
rlabel metal2 s 10314 22714 10422 22790 4 gnd
port 541 nsew
rlabel metal2 s 19050 21450 19158 21526 4 gnd
port 541 nsew
rlabel metal2 s 7050 7704 7158 7780 4 gnd
port 541 nsew
rlabel metal2 s 12042 5334 12150 5410 4 gnd
port 541 nsew
rlabel metal2 s 810 8240 918 8350 4 gnd
port 541 nsew
rlabel metal2 s 1578 1130 1686 1240 4 gnd
port 541 nsew
rlabel metal2 s 12042 14560 12150 14670 4 gnd
port 541 nsew
rlabel metal2 s 19530 3280 19638 3356 4 gnd
port 541 nsew
rlabel metal2 s 330 4544 438 4620 4 gnd
port 541 nsew
rlabel metal2 s 17802 17184 17910 17260 4 gnd
port 541 nsew
rlabel metal2 s 19050 2174 19158 2250 4 gnd
port 541 nsew
rlabel metal2 s 4554 7230 4662 7306 4 gnd
port 541 nsew
rlabel metal2 s 4074 20880 4182 20990 4 gnd
port 541 nsew
rlabel metal2 s 20778 24830 20886 24940 4 gnd
port 541 nsew
rlabel metal2 s 7050 23250 7158 23360 4 gnd
port 541 nsew
rlabel metal2 s 330 1700 438 1776 4 gnd
port 541 nsew
rlabel metal2 s 15786 594 15894 670 4 gnd
port 541 nsew
rlabel metal2 s 5322 340 5430 450 4 gnd
port 541 nsew
rlabel metal2 s 10794 23030 10902 23106 4 gnd
port 541 nsew
rlabel metal2 s 17034 15920 17142 15996 4 gnd
port 541 nsew
rlabel metal2 s 6570 2964 6678 3040 4 gnd
port 541 nsew
rlabel metal2 s 13290 6914 13398 6990 4 gnd
port 541 nsew
rlabel metal2 s 17034 20660 17142 20736 4 gnd
port 541 nsew
rlabel metal2 s 10314 10864 10422 10940 4 gnd
port 541 nsew
rlabel metal2 s 2058 3280 2166 3356 4 gnd
port 541 nsew
rlabel metal2 s 18282 18290 18390 18366 4 gnd
port 541 nsew
rlabel metal2 s 330 21924 438 22000 4 gnd
port 541 nsew
rlabel metal2 s 15306 7450 15414 7560 4 gnd
port 541 nsew
rlabel metal2 s 18282 21450 18390 21526 4 gnd
port 541 nsew
rlabel metal2 s 15786 7230 15894 7306 4 gnd
port 541 nsew
rlabel metal2 s 10314 17184 10422 17260 4 gnd
port 541 nsew
rlabel metal2 s 19050 2710 19158 2820 4 gnd
port 541 nsew
rlabel metal2 s 11562 18290 11670 18366 4 gnd
port 541 nsew
rlabel metal2 s 12810 8494 12918 8570 4 gnd
port 541 nsew
rlabel metal2 s 12042 24294 12150 24370 4 gnd
port 541 nsew
rlabel metal2 s 5802 594 5910 670 4 gnd
port 541 nsew
rlabel metal2 s 810 17184 918 17260 4 gnd
port 541 nsew
rlabel metal2 s 17802 6660 17910 6770 4 gnd
port 541 nsew
rlabel metal2 s 810 4070 918 4146 4 gnd
port 541 nsew
rlabel metal2 s 330 3500 438 3610 4 gnd
port 541 nsew
rlabel metal2 s 9066 13770 9174 13880 4 gnd
port 541 nsew
rlabel metal2 s 5802 2964 5910 3040 4 gnd
port 541 nsew
rlabel metal2 s 17802 17974 17910 18050 4 gnd
port 541 nsew
rlabel metal2 s 9066 1384 9174 1460 4 gnd
port 541 nsew
rlabel metal2 s 14058 9820 14166 9930 4 gnd
port 541 nsew
rlabel metal2 s 16554 17974 16662 18050 4 gnd
port 541 nsew
rlabel metal2 s 4554 24040 4662 24150 4 gnd
port 541 nsew
rlabel metal2 s 11562 4290 11670 4400 4 gnd
port 541 nsew
rlabel metal2 s 11562 11970 11670 12046 4 gnd
port 541 nsew
rlabel metal2 s 12810 16930 12918 17040 4 gnd
port 541 nsew
rlabel metal2 s 4074 8810 4182 8886 4 gnd
port 541 nsew
rlabel metal2 s 20298 12760 20406 12836 4 gnd
port 541 nsew
rlabel metal2 s 4074 5870 4182 5980 4 gnd
port 541 nsew
rlabel metal2 s 19530 4070 19638 4146 4 gnd
port 541 nsew
rlabel metal2 s 14538 9820 14646 9930 4 gnd
port 541 nsew
rlabel metal2 s 2826 16394 2934 16470 4 gnd
port 541 nsew
rlabel metal2 s 20298 4290 20406 4400 4 gnd
port 541 nsew
rlabel metal2 s 18282 15350 18390 15460 4 gnd
port 541 nsew
rlabel metal2 s 12042 3754 12150 3830 4 gnd
port 541 nsew
rlabel metal2 s 12042 1920 12150 2030 4 gnd
port 541 nsew
rlabel metal2 s 15306 15130 15414 15206 4 gnd
port 541 nsew
rlabel metal2 s 9546 19870 9654 19946 4 gnd
port 541 nsew
rlabel metal2 s 13290 8494 13398 8570 4 gnd
port 541 nsew
rlabel metal2 s 6570 9600 6678 9676 4 gnd
port 541 nsew
rlabel metal2 s 7050 25084 7158 25160 4 gnd
port 541 nsew
rlabel metal2 s 2058 14814 2166 14890 4 gnd
port 541 nsew
rlabel metal2 s 15306 1920 15414 2030 4 gnd
port 541 nsew
rlabel metal2 s 2826 10864 2934 10940 4 gnd
port 541 nsew
rlabel metal2 s 19050 13234 19158 13310 4 gnd
port 541 nsew
rlabel metal2 s 7050 13550 7158 13626 4 gnd
port 541 nsew
rlabel metal2 s 14058 2710 14166 2820 4 gnd
port 541 nsew
rlabel metal2 s 14538 12760 14646 12836 4 gnd
port 541 nsew
rlabel metal2 s 20778 16930 20886 17040 4 gnd
port 541 nsew
rlabel metal2 s 5802 7450 5910 7560 4 gnd
port 541 nsew
rlabel metal2 s 20298 25874 20406 25950 4 gnd
port 541 nsew
rlabel metal2 s 810 14814 918 14890 4 gnd
port 541 nsew
rlabel metal2 s 12042 16140 12150 16250 4 gnd
port 541 nsew
rlabel metal2 s 13290 15920 13398 15996 4 gnd
port 541 nsew
rlabel metal2 s 4554 17184 4662 17260 4 gnd
port 541 nsew
rlabel metal2 s 810 24294 918 24370 4 gnd
port 541 nsew
rlabel metal2 s 810 4860 918 4936 4 gnd
port 541 nsew
rlabel metal2 s 330 7704 438 7780 4 gnd
port 541 nsew
rlabel metal2 s 2826 13234 2934 13310 4 gnd
port 541 nsew
rlabel metal2 s 2826 16710 2934 16786 4 gnd
port 541 nsew
rlabel metal2 s 8298 13770 8406 13880 4 gnd
port 541 nsew
rlabel metal2 s 11562 120 11670 196 4 gnd
port 541 nsew
rlabel metal2 s 15786 16140 15894 16250 4 gnd
port 541 nsew
rlabel metal2 s 17802 16140 17910 16250 4 gnd
port 541 nsew
rlabel metal2 s 9066 8240 9174 8350 4 gnd
port 541 nsew
rlabel metal2 s 1578 17184 1686 17260 4 gnd
port 541 nsew
rlabel metal2 s 20298 24294 20406 24370 4 gnd
port 541 nsew
rlabel metal2 s 4554 21670 4662 21780 4 gnd
port 541 nsew
rlabel metal2 s 15306 14560 15414 14670 4 gnd
port 541 nsew
rlabel metal2 s 1578 17500 1686 17576 4 gnd
port 541 nsew
rlabel metal2 s 19050 16394 19158 16470 4 gnd
port 541 nsew
rlabel metal2 s 7050 7450 7158 7560 4 gnd
port 541 nsew
rlabel metal2 s 14538 13234 14646 13310 4 gnd
port 541 nsew
rlabel metal2 s 9546 4290 9654 4400 4 gnd
port 541 nsew
rlabel metal2 s 19530 15604 19638 15680 4 gnd
port 541 nsew
rlabel metal2 s 330 23030 438 23106 4 gnd
port 541 nsew
rlabel metal2 s 12042 4860 12150 4936 4 gnd
port 541 nsew
rlabel metal2 s 12810 10610 12918 10720 4 gnd
port 541 nsew
rlabel metal2 s 17034 8810 17142 8886 4 gnd
port 541 nsew
rlabel metal2 s 20298 5334 20406 5410 4 gnd
port 541 nsew
rlabel metal2 s 1578 8810 1686 8886 4 gnd
port 541 nsew
rlabel metal2 s 17034 21134 17142 21210 4 gnd
port 541 nsew
rlabel metal2 s 9546 24040 9654 24150 4 gnd
port 541 nsew
rlabel metal2 s 20298 594 20406 670 4 gnd
port 541 nsew
rlabel metal2 s 17802 3500 17910 3610 4 gnd
port 541 nsew
rlabel metal2 s 7050 21670 7158 21780 4 gnd
port 541 nsew
rlabel metal2 s 7050 1130 7158 1240 4 gnd
port 541 nsew
rlabel metal2 s 8298 11970 8406 12046 4 gnd
port 541 nsew
rlabel metal2 s 14058 7230 14166 7306 4 gnd
port 541 nsew
rlabel metal2 s 1578 20660 1686 20736 4 gnd
port 541 nsew
rlabel metal2 s 20778 14560 20886 14670 4 gnd
port 541 nsew
rlabel metal2 s 330 16710 438 16786 4 gnd
port 541 nsew
rlabel metal2 s 10314 13234 10422 13310 4 gnd
port 541 nsew
rlabel metal2 s 8298 6660 8406 6770 4 gnd
port 541 nsew
rlabel metal2 s 19530 6914 19638 6990 4 gnd
port 541 nsew
rlabel metal2 s 12042 16930 12150 17040 4 gnd
port 541 nsew
rlabel metal2 s 15786 12760 15894 12836 4 gnd
port 541 nsew
rlabel metal2 s 1578 14340 1686 14416 4 gnd
port 541 nsew
rlabel metal2 s 20778 4860 20886 4936 4 gnd
port 541 nsew
rlabel metal2 s 9546 7230 9654 7306 4 gnd
port 541 nsew
rlabel metal2 s 2826 9600 2934 9676 4 gnd
port 541 nsew
rlabel metal2 s 16554 23250 16662 23360 4 gnd
port 541 nsew
rlabel metal2 s 16554 22714 16662 22790 4 gnd
port 541 nsew
rlabel metal2 s 14058 8494 14166 8570 4 gnd
port 541 nsew
rlabel metal2 s 2826 19300 2934 19410 4 gnd
port 541 nsew
rlabel metal2 s 10314 25620 10422 25730 4 gnd
port 541 nsew
rlabel metal2 s 810 12760 918 12836 4 gnd
port 541 nsew
rlabel metal2 s 17034 10864 17142 10940 4 gnd
port 541 nsew
rlabel metal2 s 15786 9820 15894 9930 4 gnd
port 541 nsew
rlabel metal2 s 12810 3280 12918 3356 4 gnd
port 541 nsew
rlabel metal2 s 19050 11970 19158 12046 4 gnd
port 541 nsew
rlabel metal2 s 2826 340 2934 450 4 gnd
port 541 nsew
rlabel metal2 s 9066 24040 9174 24150 4 gnd
port 541 nsew
rlabel metal2 s 15786 15130 15894 15206 4 gnd
port 541 nsew
rlabel metal2 s 17034 18764 17142 18840 4 gnd
port 541 nsew
rlabel metal2 s 7050 23504 7158 23580 4 gnd
port 541 nsew
rlabel metal2 s 7818 4860 7926 4936 4 gnd
port 541 nsew
rlabel metal2 s 6570 23030 6678 23106 4 gnd
port 541 nsew
rlabel metal2 s 2058 19554 2166 19630 4 gnd
port 541 nsew
rlabel metal2 s 810 22240 918 22316 4 gnd
port 541 nsew
rlabel metal2 s 15786 6914 15894 6990 4 gnd
port 541 nsew
rlabel metal2 s 20778 15350 20886 15460 4 gnd
port 541 nsew
rlabel metal2 s 3306 22460 3414 22570 4 gnd
port 541 nsew
rlabel metal2 s 1578 21924 1686 22000 4 gnd
port 541 nsew
rlabel metal2 s 17034 15604 17142 15680 4 gnd
port 541 nsew
rlabel metal2 s 4554 5080 4662 5190 4 gnd
port 541 nsew
rlabel metal2 s 6570 17974 6678 18050 4 gnd
port 541 nsew
rlabel metal2 s 10794 20660 10902 20736 4 gnd
port 541 nsew
rlabel metal2 s 13290 18510 13398 18620 4 gnd
port 541 nsew
rlabel metal2 s 2826 14814 2934 14890 4 gnd
port 541 nsew
rlabel metal2 s 17034 20344 17142 20420 4 gnd
port 541 nsew
rlabel metal2 s 2058 1700 2166 1776 4 gnd
port 541 nsew
rlabel metal2 s 10794 8240 10902 8350 4 gnd
port 541 nsew
rlabel metal2 s 20298 23504 20406 23580 4 gnd
port 541 nsew
rlabel metal2 s 12042 21134 12150 21210 4 gnd
port 541 nsew
rlabel metal2 s 10794 19080 10902 19156 4 gnd
port 541 nsew
rlabel metal2 s 810 10864 918 10940 4 gnd
port 541 nsew
rlabel metal2 s 2826 9030 2934 9140 4 gnd
port 541 nsew
rlabel metal2 s 14538 2710 14646 2820 4 gnd
port 541 nsew
rlabel metal2 s 7050 20090 7158 20200 4 gnd
port 541 nsew
rlabel metal2 s 17802 8020 17910 8096 4 gnd
port 541 nsew
rlabel metal2 s 15306 10074 15414 10150 4 gnd
port 541 nsew
rlabel metal2 s 1578 12190 1686 12300 4 gnd
port 541 nsew
rlabel metal2 s 8298 3500 8406 3610 4 gnd
port 541 nsew
rlabel metal2 s 14538 21134 14646 21210 4 gnd
port 541 nsew
rlabel metal2 s 8298 25874 8406 25950 4 gnd
port 541 nsew
rlabel metal2 s 5322 22714 5430 22790 4 gnd
port 541 nsew
rlabel metal2 s 2826 17974 2934 18050 4 gnd
port 541 nsew
rlabel metal2 s 3306 3280 3414 3356 4 gnd
port 541 nsew
rlabel metal2 s 3306 18764 3414 18840 4 gnd
port 541 nsew
rlabel metal2 s 6570 14560 6678 14670 4 gnd
port 541 nsew
rlabel metal2 s 2826 3280 2934 3356 4 gnd
port 541 nsew
rlabel metal2 s 15786 24610 15894 24686 4 gnd
port 541 nsew
rlabel metal2 s 330 594 438 670 4 gnd
port 541 nsew
rlabel metal2 s 12810 13550 12918 13626 4 gnd
port 541 nsew
rlabel metal2 s 330 11400 438 11510 4 gnd
port 541 nsew
rlabel metal2 s 10794 21450 10902 21526 4 gnd
port 541 nsew
rlabel metal2 s 4554 17720 4662 17830 4 gnd
port 541 nsew
rlabel metal2 s 810 23030 918 23106 4 gnd
port 541 nsew
rlabel metal2 s 10314 25084 10422 25160 4 gnd
port 541 nsew
rlabel metal2 s 18282 5080 18390 5190 4 gnd
port 541 nsew
rlabel metal2 s 5322 4070 5430 4146 4 gnd
port 541 nsew
rlabel metal2 s 14538 23030 14646 23106 4 gnd
port 541 nsew
rlabel metal2 s 20298 10864 20406 10940 4 gnd
port 541 nsew
rlabel metal2 s 16554 2174 16662 2250 4 gnd
port 541 nsew
rlabel metal2 s 8298 23030 8406 23106 4 gnd
port 541 nsew
rlabel metal2 s 6570 11654 6678 11730 4 gnd
port 541 nsew
rlabel metal2 s 7818 7450 7926 7560 4 gnd
port 541 nsew
rlabel metal2 s 18282 18764 18390 18840 4 gnd
port 541 nsew
rlabel metal2 s 20778 9600 20886 9676 4 gnd
port 541 nsew
rlabel metal2 s 9546 7450 9654 7560 4 gnd
port 541 nsew
rlabel metal2 s 12042 9820 12150 9930 4 gnd
port 541 nsew
rlabel metal2 s 9066 21670 9174 21780 4 gnd
port 541 nsew
rlabel metal2 s 15786 23030 15894 23106 4 gnd
port 541 nsew
rlabel metal2 s 13290 3754 13398 3830 4 gnd
port 541 nsew
rlabel metal2 s 9546 12980 9654 13090 4 gnd
port 541 nsew
rlabel metal2 s 19530 20660 19638 20736 4 gnd
port 541 nsew
rlabel metal2 s 20298 7704 20406 7780 4 gnd
port 541 nsew
rlabel metal2 s 3306 15920 3414 15996 4 gnd
port 541 nsew
rlabel metal2 s 12810 6124 12918 6200 4 gnd
port 541 nsew
rlabel metal2 s 4554 15350 4662 15460 4 gnd
port 541 nsew
rlabel metal2 s 13290 4860 13398 4936 4 gnd
port 541 nsew
rlabel metal2 s 4554 594 4662 670 4 gnd
port 541 nsew
rlabel metal2 s 1578 17720 1686 17830 4 gnd
port 541 nsew
rlabel metal2 s 5802 23504 5910 23580 4 gnd
port 541 nsew
rlabel metal2 s 13290 22714 13398 22790 4 gnd
port 541 nsew
rlabel metal2 s 6570 25400 6678 25476 4 gnd
port 541 nsew
rlabel metal2 s 11562 3500 11670 3610 4 gnd
port 541 nsew
rlabel metal2 s 10314 18764 10422 18840 4 gnd
port 541 nsew
rlabel metal2 s 19530 9030 19638 9140 4 gnd
port 541 nsew
rlabel metal2 s 8298 21134 8406 21210 4 gnd
port 541 nsew
rlabel metal2 s 2826 4070 2934 4146 4 gnd
port 541 nsew
rlabel metal2 s 12042 1384 12150 1460 4 gnd
port 541 nsew
rlabel metal2 s 3306 21670 3414 21780 4 gnd
port 541 nsew
rlabel metal2 s 20778 16710 20886 16786 4 gnd
port 541 nsew
rlabel metal2 s 11562 7450 11670 7560 4 gnd
port 541 nsew
rlabel metal2 s 330 9600 438 9676 4 gnd
port 541 nsew
rlabel metal2 s 12810 18764 12918 18840 4 gnd
port 541 nsew
rlabel metal2 s 14538 18290 14646 18366 4 gnd
port 541 nsew
rlabel metal2 s 20298 3280 20406 3356 4 gnd
port 541 nsew
rlabel metal2 s 12810 4544 12918 4620 4 gnd
port 541 nsew
rlabel metal2 s 13290 4544 13398 4620 4 gnd
port 541 nsew
rlabel metal2 s 4554 15130 4662 15206 4 gnd
port 541 nsew
rlabel metal2 s 6570 24294 6678 24370 4 gnd
port 541 nsew
rlabel metal2 s 9546 2490 9654 2566 4 gnd
port 541 nsew
rlabel metal2 s 5322 2174 5430 2250 4 gnd
port 541 nsew
rlabel metal2 s 810 1130 918 1240 4 gnd
port 541 nsew
rlabel metal2 s 7818 4290 7926 4400 4 gnd
port 541 nsew
rlabel metal2 s 15306 4860 15414 4936 4 gnd
port 541 nsew
rlabel metal2 s 10794 4860 10902 4936 4 gnd
port 541 nsew
rlabel metal2 s 19050 18764 19158 18840 4 gnd
port 541 nsew
rlabel metal2 s 10794 24830 10902 24940 4 gnd
port 541 nsew
rlabel metal2 s 1578 2710 1686 2820 4 gnd
port 541 nsew
rlabel metal2 s 10794 15604 10902 15680 4 gnd
port 541 nsew
rlabel metal2 s 16554 8494 16662 8570 4 gnd
port 541 nsew
rlabel metal2 s 9546 3754 9654 3830 4 gnd
port 541 nsew
rlabel metal2 s 20778 23250 20886 23360 4 gnd
port 541 nsew
rlabel metal2 s 13290 2710 13398 2820 4 gnd
port 541 nsew
rlabel metal2 s 11562 17500 11670 17576 4 gnd
port 541 nsew
rlabel metal2 s 9066 25084 9174 25160 4 gnd
port 541 nsew
rlabel metal2 s 3306 3754 3414 3830 4 gnd
port 541 nsew
rlabel metal2 s 12810 24294 12918 24370 4 gnd
port 541 nsew
rlabel metal2 s 9546 10390 9654 10466 4 gnd
port 541 nsew
rlabel metal2 s 2826 20090 2934 20200 4 gnd
port 541 nsew
rlabel metal2 s 15306 24610 15414 24686 4 gnd
port 541 nsew
rlabel metal2 s 17034 2490 17142 2566 4 gnd
port 541 nsew
rlabel metal2 s 18282 5650 18390 5726 4 gnd
port 541 nsew
rlabel metal2 s 2826 5080 2934 5190 4 gnd
port 541 nsew
rlabel metal2 s 5802 20090 5910 20200 4 gnd
port 541 nsew
rlabel metal2 s 16554 23030 16662 23106 4 gnd
port 541 nsew
rlabel metal2 s 9546 12760 9654 12836 4 gnd
port 541 nsew
rlabel metal2 s 8298 12980 8406 13090 4 gnd
port 541 nsew
rlabel metal2 s 9066 594 9174 670 4 gnd
port 541 nsew
rlabel metal2 s 14058 18290 14166 18366 4 gnd
port 541 nsew
rlabel metal2 s 7818 18764 7926 18840 4 gnd
port 541 nsew
rlabel metal2 s 16554 15604 16662 15680 4 gnd
port 541 nsew
rlabel metal2 s 1578 16394 1686 16470 4 gnd
port 541 nsew
rlabel metal2 s 17802 19554 17910 19630 4 gnd
port 541 nsew
rlabel metal2 s 6570 11180 6678 11256 4 gnd
port 541 nsew
rlabel metal2 s 18282 594 18390 670 4 gnd
port 541 nsew
rlabel metal2 s 330 24294 438 24370 4 gnd
port 541 nsew
rlabel metal2 s 2058 10864 2166 10940 4 gnd
port 541 nsew
rlabel metal2 s 4554 20090 4662 20200 4 gnd
port 541 nsew
rlabel metal2 s 330 6440 438 6516 4 gnd
port 541 nsew
rlabel metal2 s 20298 5080 20406 5190 4 gnd
port 541 nsew
rlabel metal2 s 20298 6914 20406 6990 4 gnd
port 541 nsew
rlabel metal2 s 19530 4544 19638 4620 4 gnd
port 541 nsew
rlabel metal2 s 16554 11970 16662 12046 4 gnd
port 541 nsew
rlabel metal2 s 10794 16394 10902 16470 4 gnd
port 541 nsew
rlabel metal2 s 2826 1130 2934 1240 4 gnd
port 541 nsew
rlabel metal2 s 19530 7450 19638 7560 4 gnd
port 541 nsew
rlabel metal2 s 11562 18510 11670 18620 4 gnd
port 541 nsew
rlabel metal2 s 4554 6660 4662 6770 4 gnd
port 541 nsew
rlabel metal2 s 5802 21670 5910 21780 4 gnd
port 541 nsew
rlabel metal2 s 2826 21924 2934 22000 4 gnd
port 541 nsew
rlabel metal2 s 12042 594 12150 670 4 gnd
port 541 nsew
rlabel metal2 s 6570 21450 6678 21526 4 gnd
port 541 nsew
rlabel metal2 s 17034 12980 17142 13090 4 gnd
port 541 nsew
rlabel metal2 s 19050 16710 19158 16786 4 gnd
port 541 nsew
rlabel metal2 s 19050 23250 19158 23360 4 gnd
port 541 nsew
rlabel metal2 s 16554 14560 16662 14670 4 gnd
port 541 nsew
rlabel metal2 s 7050 5334 7158 5410 4 gnd
port 541 nsew
rlabel metal2 s 4074 9030 4182 9140 4 gnd
port 541 nsew
rlabel metal2 s 3306 15604 3414 15680 4 gnd
port 541 nsew
rlabel metal2 s 4554 17500 4662 17576 4 gnd
port 541 nsew
rlabel metal2 s 14058 22714 14166 22790 4 gnd
port 541 nsew
rlabel metal2 s 1578 20090 1686 20200 4 gnd
port 541 nsew
rlabel metal2 s 12810 5080 12918 5190 4 gnd
port 541 nsew
rlabel metal2 s 14058 25084 14166 25160 4 gnd
port 541 nsew
rlabel metal2 s 2058 24040 2166 24150 4 gnd
port 541 nsew
rlabel metal2 s 10794 25620 10902 25730 4 gnd
port 541 nsew
rlabel metal2 s 19050 10074 19158 10150 4 gnd
port 541 nsew
rlabel metal2 s 9066 16930 9174 17040 4 gnd
port 541 nsew
rlabel metal2 s 14538 14814 14646 14890 4 gnd
port 541 nsew
rlabel metal2 s 8298 22714 8406 22790 4 gnd
port 541 nsew
rlabel metal2 s 10314 16394 10422 16470 4 gnd
port 541 nsew
rlabel metal2 s 19530 15350 19638 15460 4 gnd
port 541 nsew
rlabel metal2 s 18282 6914 18390 6990 4 gnd
port 541 nsew
rlabel metal2 s 7050 4860 7158 4936 4 gnd
port 541 nsew
rlabel metal2 s 12810 9284 12918 9360 4 gnd
port 541 nsew
rlabel metal2 s 4074 11654 4182 11730 4 gnd
port 541 nsew
rlabel metal2 s 15786 1384 15894 1460 4 gnd
port 541 nsew
rlabel metal2 s 18282 21134 18390 21210 4 gnd
port 541 nsew
rlabel metal2 s 17034 1920 17142 2030 4 gnd
port 541 nsew
rlabel metal2 s 1578 1920 1686 2030 4 gnd
port 541 nsew
rlabel metal2 s 7818 24830 7926 24940 4 gnd
port 541 nsew
rlabel metal2 s 19050 5870 19158 5980 4 gnd
port 541 nsew
rlabel metal2 s 12042 21450 12150 21526 4 gnd
port 541 nsew
rlabel metal2 s 11562 23250 11670 23360 4 gnd
port 541 nsew
rlabel metal2 s 18282 3754 18390 3830 4 gnd
port 541 nsew
rlabel metal2 s 330 13770 438 13880 4 gnd
port 541 nsew
rlabel metal2 s 17802 12190 17910 12300 4 gnd
port 541 nsew
rlabel metal2 s 10794 20880 10902 20990 4 gnd
port 541 nsew
rlabel metal2 s 16554 21924 16662 22000 4 gnd
port 541 nsew
rlabel metal2 s 8298 9284 8406 9360 4 gnd
port 541 nsew
rlabel metal2 s 330 14814 438 14890 4 gnd
port 541 nsew
rlabel metal2 s 20778 3754 20886 3830 4 gnd
port 541 nsew
rlabel metal2 s 8298 8810 8406 8886 4 gnd
port 541 nsew
rlabel metal2 s 14058 5334 14166 5410 4 gnd
port 541 nsew
rlabel metal2 s 17802 21134 17910 21210 4 gnd
port 541 nsew
rlabel metal2 s 2058 6124 2166 6200 4 gnd
port 541 nsew
rlabel metal2 s 9066 12980 9174 13090 4 gnd
port 541 nsew
rlabel metal2 s 9546 18510 9654 18620 4 gnd
port 541 nsew
rlabel metal2 s 20298 8020 20406 8096 4 gnd
port 541 nsew
rlabel metal2 s 4554 25620 4662 25730 4 gnd
port 541 nsew
rlabel metal2 s 6570 12980 6678 13090 4 gnd
port 541 nsew
rlabel metal2 s 15786 15604 15894 15680 4 gnd
port 541 nsew
rlabel metal2 s 10794 120 10902 196 4 gnd
port 541 nsew
rlabel metal2 s 4554 4860 4662 4936 4 gnd
port 541 nsew
rlabel metal2 s 19530 17500 19638 17576 4 gnd
port 541 nsew
rlabel metal2 s 17034 16394 17142 16470 4 gnd
port 541 nsew
rlabel metal2 s 9066 6660 9174 6770 4 gnd
port 541 nsew
rlabel metal2 s 9546 14814 9654 14890 4 gnd
port 541 nsew
rlabel metal2 s 14538 15350 14646 15460 4 gnd
port 541 nsew
rlabel metal2 s 15786 22240 15894 22316 4 gnd
port 541 nsew
rlabel metal2 s 8298 9600 8406 9676 4 gnd
port 541 nsew
rlabel metal2 s 10794 8020 10902 8096 4 gnd
port 541 nsew
rlabel metal2 s 10314 3754 10422 3830 4 gnd
port 541 nsew
rlabel metal2 s 19050 120 19158 196 4 gnd
port 541 nsew
rlabel metal2 s 20298 20344 20406 20420 4 gnd
port 541 nsew
rlabel metal2 s 2058 17184 2166 17260 4 gnd
port 541 nsew
rlabel metal2 s 7818 15130 7926 15206 4 gnd
port 541 nsew
rlabel metal2 s 13290 19080 13398 19156 4 gnd
port 541 nsew
rlabel metal2 s 20298 14340 20406 14416 4 gnd
port 541 nsew
rlabel metal2 s 4554 5870 4662 5980 4 gnd
port 541 nsew
rlabel metal2 s 8298 5650 8406 5726 4 gnd
port 541 nsew
rlabel metal2 s 15306 16394 15414 16470 4 gnd
port 541 nsew
rlabel metal2 s 8298 3754 8406 3830 4 gnd
port 541 nsew
rlabel metal2 s 330 3754 438 3830 4 gnd
port 541 nsew
rlabel metal2 s 17034 25620 17142 25730 4 gnd
port 541 nsew
rlabel metal2 s 18282 14340 18390 14416 4 gnd
port 541 nsew
rlabel metal2 s 19530 120 19638 196 4 gnd
port 541 nsew
rlabel metal2 s 2058 4290 2166 4400 4 gnd
port 541 nsew
rlabel metal2 s 3306 594 3414 670 4 gnd
port 541 nsew
rlabel metal2 s 17802 17500 17910 17576 4 gnd
port 541 nsew
rlabel metal2 s 3306 22240 3414 22316 4 gnd
port 541 nsew
rlabel metal2 s 2826 6914 2934 6990 4 gnd
port 541 nsew
rlabel metal2 s 4074 10610 4182 10720 4 gnd
port 541 nsew
rlabel metal2 s 19530 3500 19638 3610 4 gnd
port 541 nsew
rlabel metal2 s 8298 17184 8406 17260 4 gnd
port 541 nsew
rlabel metal2 s 330 15920 438 15996 4 gnd
port 541 nsew
rlabel metal2 s 12042 25874 12150 25950 4 gnd
port 541 nsew
rlabel metal2 s 20298 24040 20406 24150 4 gnd
port 541 nsew
rlabel metal2 s 1578 23504 1686 23580 4 gnd
port 541 nsew
rlabel metal2 s 15306 5650 15414 5726 4 gnd
port 541 nsew
rlabel metal2 s 8298 8020 8406 8096 4 gnd
port 541 nsew
rlabel metal2 s 2826 17500 2934 17576 4 gnd
port 541 nsew
rlabel metal2 s 6570 25874 6678 25950 4 gnd
port 541 nsew
rlabel metal2 s 4074 21134 4182 21210 4 gnd
port 541 nsew
rlabel metal2 s 9546 22240 9654 22316 4 gnd
port 541 nsew
rlabel metal2 s 19050 5650 19158 5726 4 gnd
port 541 nsew
rlabel metal2 s 17802 21450 17910 21526 4 gnd
port 541 nsew
rlabel metal2 s 12810 5870 12918 5980 4 gnd
port 541 nsew
rlabel metal2 s 810 11180 918 11256 4 gnd
port 541 nsew
rlabel metal2 s 8298 14814 8406 14890 4 gnd
port 541 nsew
rlabel metal2 s 18282 24830 18390 24940 4 gnd
port 541 nsew
rlabel metal2 s 11562 17184 11670 17260 4 gnd
port 541 nsew
rlabel metal2 s 12042 16710 12150 16786 4 gnd
port 541 nsew
rlabel metal2 s 5802 21134 5910 21210 4 gnd
port 541 nsew
rlabel metal2 s 7050 3280 7158 3356 4 gnd
port 541 nsew
rlabel metal2 s 19530 14814 19638 14890 4 gnd
port 541 nsew
rlabel metal2 s 15306 19080 15414 19156 4 gnd
port 541 nsew
rlabel metal2 s 18282 340 18390 450 4 gnd
port 541 nsew
rlabel metal2 s 3306 1384 3414 1460 4 gnd
port 541 nsew
rlabel metal2 s 18282 22714 18390 22790 4 gnd
port 541 nsew
rlabel metal2 s 10794 25874 10902 25950 4 gnd
port 541 nsew
rlabel metal2 s 810 8020 918 8096 4 gnd
port 541 nsew
rlabel metal2 s 18282 5334 18390 5410 4 gnd
port 541 nsew
rlabel metal2 s 5802 12190 5910 12300 4 gnd
port 541 nsew
rlabel metal2 s 15306 9820 15414 9930 4 gnd
port 541 nsew
rlabel metal2 s 19530 1130 19638 1240 4 gnd
port 541 nsew
rlabel metal2 s 20778 25400 20886 25476 4 gnd
port 541 nsew
rlabel metal2 s 810 6914 918 6990 4 gnd
port 541 nsew
rlabel metal2 s 12810 9600 12918 9676 4 gnd
port 541 nsew
rlabel metal2 s 5322 1384 5430 1460 4 gnd
port 541 nsew
rlabel metal2 s 15786 5870 15894 5980 4 gnd
port 541 nsew
rlabel metal2 s 4074 17720 4182 17830 4 gnd
port 541 nsew
rlabel metal2 s 20298 21670 20406 21780 4 gnd
port 541 nsew
rlabel metal2 s 2058 22240 2166 22316 4 gnd
port 541 nsew
rlabel metal2 s 20298 4070 20406 4146 4 gnd
port 541 nsew
rlabel metal2 s 9066 11654 9174 11730 4 gnd
port 541 nsew
rlabel metal2 s 5322 17974 5430 18050 4 gnd
port 541 nsew
rlabel metal2 s 14058 12444 14166 12520 4 gnd
port 541 nsew
rlabel metal2 s 6570 8810 6678 8886 4 gnd
port 541 nsew
rlabel metal2 s 12042 11400 12150 11510 4 gnd
port 541 nsew
rlabel metal2 s 1578 21450 1686 21526 4 gnd
port 541 nsew
rlabel metal2 s 10314 9030 10422 9140 4 gnd
port 541 nsew
rlabel metal2 s 1578 18290 1686 18366 4 gnd
port 541 nsew
rlabel metal2 s 15786 3500 15894 3610 4 gnd
port 541 nsew
rlabel metal2 s 20298 11654 20406 11730 4 gnd
port 541 nsew
rlabel metal2 s 7050 2174 7158 2250 4 gnd
port 541 nsew
rlabel metal2 s 4074 19554 4182 19630 4 gnd
port 541 nsew
rlabel metal2 s 18282 7704 18390 7780 4 gnd
port 541 nsew
rlabel metal2 s 15786 17720 15894 17830 4 gnd
port 541 nsew
rlabel metal2 s 10794 19554 10902 19630 4 gnd
port 541 nsew
rlabel metal2 s 6570 5870 6678 5980 4 gnd
port 541 nsew
rlabel metal2 s 10314 11970 10422 12046 4 gnd
port 541 nsew
rlabel metal2 s 4074 7450 4182 7560 4 gnd
port 541 nsew
rlabel metal2 s 2058 2490 2166 2566 4 gnd
port 541 nsew
rlabel metal2 s 12042 25084 12150 25160 4 gnd
port 541 nsew
rlabel metal2 s 5802 23250 5910 23360 4 gnd
port 541 nsew
rlabel metal2 s 1578 5870 1686 5980 4 gnd
port 541 nsew
rlabel metal2 s 13290 2964 13398 3040 4 gnd
port 541 nsew
rlabel metal2 s 17802 7450 17910 7560 4 gnd
port 541 nsew
rlabel metal2 s 6570 1384 6678 1460 4 gnd
port 541 nsew
rlabel metal2 s 14538 19300 14646 19410 4 gnd
port 541 nsew
rlabel metal2 s 4074 25620 4182 25730 4 gnd
port 541 nsew
rlabel metal2 s 20298 15350 20406 15460 4 gnd
port 541 nsew
rlabel metal2 s 1578 15350 1686 15460 4 gnd
port 541 nsew
rlabel metal2 s 5322 4544 5430 4620 4 gnd
port 541 nsew
rlabel metal2 s 10794 2710 10902 2820 4 gnd
port 541 nsew
rlabel metal2 s 15306 25084 15414 25160 4 gnd
port 541 nsew
rlabel metal2 s 20298 24610 20406 24686 4 gnd
port 541 nsew
rlabel metal2 s 12042 14340 12150 14416 4 gnd
port 541 nsew
rlabel metal2 s 20298 11180 20406 11256 4 gnd
port 541 nsew
rlabel metal2 s 20778 7704 20886 7780 4 gnd
port 541 nsew
rlabel metal2 s 13290 5650 13398 5726 4 gnd
port 541 nsew
rlabel metal2 s 1578 21134 1686 21210 4 gnd
port 541 nsew
rlabel metal2 s 3306 17184 3414 17260 4 gnd
port 541 nsew
rlabel metal2 s 7050 4544 7158 4620 4 gnd
port 541 nsew
rlabel metal2 s 4554 24294 4662 24370 4 gnd
port 541 nsew
rlabel metal2 s 4074 17974 4182 18050 4 gnd
port 541 nsew
rlabel metal2 s 1578 14560 1686 14670 4 gnd
port 541 nsew
rlabel metal2 s 6570 20880 6678 20990 4 gnd
port 541 nsew
rlabel metal2 s 14538 15604 14646 15680 4 gnd
port 541 nsew
rlabel metal2 s 14058 1920 14166 2030 4 gnd
port 541 nsew
rlabel metal2 s 13290 5870 13398 5980 4 gnd
port 541 nsew
rlabel metal2 s 5322 2710 5430 2820 4 gnd
port 541 nsew
rlabel metal2 s 810 16394 918 16470 4 gnd
port 541 nsew
rlabel metal2 s 9066 18764 9174 18840 4 gnd
port 541 nsew
rlabel metal2 s 10794 23504 10902 23580 4 gnd
port 541 nsew
rlabel metal2 s 7050 9284 7158 9360 4 gnd
port 541 nsew
rlabel metal2 s 8298 11180 8406 11256 4 gnd
port 541 nsew
rlabel metal2 s 2826 5334 2934 5410 4 gnd
port 541 nsew
rlabel metal2 s 6570 1130 6678 1240 4 gnd
port 541 nsew
rlabel metal2 s 2058 2710 2166 2820 4 gnd
port 541 nsew
rlabel metal2 s 5802 9284 5910 9360 4 gnd
port 541 nsew
rlabel metal2 s 18282 4290 18390 4400 4 gnd
port 541 nsew
rlabel metal2 s 13290 23250 13398 23360 4 gnd
port 541 nsew
rlabel metal2 s 9066 7230 9174 7306 4 gnd
port 541 nsew
rlabel metal2 s 16554 12190 16662 12300 4 gnd
port 541 nsew
rlabel metal2 s 3306 19080 3414 19156 4 gnd
port 541 nsew
rlabel metal2 s 17802 9284 17910 9360 4 gnd
port 541 nsew
rlabel metal2 s 14538 18510 14646 18620 4 gnd
port 541 nsew
rlabel metal2 s 4074 6124 4182 6200 4 gnd
port 541 nsew
rlabel metal2 s 3306 17720 3414 17830 4 gnd
port 541 nsew
rlabel metal2 s 5802 16394 5910 16470 4 gnd
port 541 nsew
rlabel metal2 s 17034 9284 17142 9360 4 gnd
port 541 nsew
rlabel metal2 s 7818 20660 7926 20736 4 gnd
port 541 nsew
rlabel metal2 s 20778 6660 20886 6770 4 gnd
port 541 nsew
rlabel metal2 s 4554 4290 4662 4400 4 gnd
port 541 nsew
rlabel metal2 s 2058 16140 2166 16250 4 gnd
port 541 nsew
rlabel metal2 s 3306 5650 3414 5726 4 gnd
port 541 nsew
rlabel metal2 s 12810 4860 12918 4936 4 gnd
port 541 nsew
rlabel metal2 s 12810 24830 12918 24940 4 gnd
port 541 nsew
rlabel metal2 s 10314 20090 10422 20200 4 gnd
port 541 nsew
rlabel metal2 s 6570 14024 6678 14100 4 gnd
port 541 nsew
rlabel metal2 s 17034 3280 17142 3356 4 gnd
port 541 nsew
rlabel metal2 s 3306 4290 3414 4400 4 gnd
port 541 nsew
rlabel metal2 s 19050 25620 19158 25730 4 gnd
port 541 nsew
rlabel metal2 s 4554 3754 4662 3830 4 gnd
port 541 nsew
rlabel metal2 s 1578 24040 1686 24150 4 gnd
port 541 nsew
rlabel metal2 s 15786 17500 15894 17576 4 gnd
port 541 nsew
rlabel metal2 s 330 5650 438 5726 4 gnd
port 541 nsew
rlabel metal2 s 8298 6124 8406 6200 4 gnd
port 541 nsew
rlabel metal2 s 13290 22240 13398 22316 4 gnd
port 541 nsew
rlabel metal2 s 2058 4544 2166 4620 4 gnd
port 541 nsew
rlabel metal2 s 6570 2490 6678 2566 4 gnd
port 541 nsew
rlabel metal2 s 20778 1700 20886 1776 4 gnd
port 541 nsew
rlabel metal2 s 14058 120 14166 196 4 gnd
port 541 nsew
rlabel metal2 s 14058 2490 14166 2566 4 gnd
port 541 nsew
rlabel metal2 s 14538 14340 14646 14416 4 gnd
port 541 nsew
rlabel metal2 s 9066 12444 9174 12520 4 gnd
port 541 nsew
rlabel metal2 s 15786 1700 15894 1776 4 gnd
port 541 nsew
rlabel metal2 s 4554 25874 4662 25950 4 gnd
port 541 nsew
rlabel metal2 s 4554 20660 4662 20736 4 gnd
port 541 nsew
rlabel metal2 s 7818 25620 7926 25730 4 gnd
port 541 nsew
rlabel metal2 s 9546 23250 9654 23360 4 gnd
port 541 nsew
rlabel metal2 s 4554 16394 4662 16470 4 gnd
port 541 nsew
rlabel metal2 s 17802 11180 17910 11256 4 gnd
port 541 nsew
rlabel metal2 s 9066 22714 9174 22790 4 gnd
port 541 nsew
rlabel metal2 s 10314 18290 10422 18366 4 gnd
port 541 nsew
rlabel metal2 s 20298 6124 20406 6200 4 gnd
port 541 nsew
rlabel metal2 s 15786 15350 15894 15460 4 gnd
port 541 nsew
rlabel metal2 s 810 910 918 986 4 gnd
port 541 nsew
rlabel metal2 s 14538 594 14646 670 4 gnd
port 541 nsew
rlabel metal2 s 19050 6914 19158 6990 4 gnd
port 541 nsew
rlabel metal2 s 5802 3280 5910 3356 4 gnd
port 541 nsew
rlabel metal2 s 17802 15604 17910 15680 4 gnd
port 541 nsew
rlabel metal2 s 15306 1700 15414 1776 4 gnd
port 541 nsew
rlabel metal2 s 12810 20344 12918 20420 4 gnd
port 541 nsew
rlabel metal2 s 7818 19080 7926 19156 4 gnd
port 541 nsew
rlabel metal2 s 5322 21134 5430 21210 4 gnd
port 541 nsew
rlabel metal2 s 13290 24294 13398 24370 4 gnd
port 541 nsew
rlabel metal2 s 20778 23030 20886 23106 4 gnd
port 541 nsew
rlabel metal2 s 2826 21134 2934 21210 4 gnd
port 541 nsew
rlabel metal2 s 11562 6440 11670 6516 4 gnd
port 541 nsew
rlabel metal2 s 330 8020 438 8096 4 gnd
port 541 nsew
rlabel metal2 s 2058 19300 2166 19410 4 gnd
port 541 nsew
rlabel metal2 s 4074 340 4182 450 4 gnd
port 541 nsew
rlabel metal2 s 1578 20880 1686 20990 4 gnd
port 541 nsew
rlabel metal2 s 20778 21924 20886 22000 4 gnd
port 541 nsew
rlabel metal2 s 7050 5080 7158 5190 4 gnd
port 541 nsew
rlabel metal2 s 13290 16930 13398 17040 4 gnd
port 541 nsew
rlabel metal2 s 10314 10390 10422 10466 4 gnd
port 541 nsew
rlabel metal2 s 9546 18290 9654 18366 4 gnd
port 541 nsew
rlabel metal2 s 19050 12190 19158 12300 4 gnd
port 541 nsew
rlabel metal2 s 20298 19300 20406 19410 4 gnd
port 541 nsew
rlabel metal2 s 15786 10390 15894 10466 4 gnd
port 541 nsew
rlabel metal2 s 18282 14024 18390 14100 4 gnd
port 541 nsew
rlabel metal2 s 10794 22240 10902 22316 4 gnd
port 541 nsew
rlabel metal2 s 4074 6914 4182 6990 4 gnd
port 541 nsew
rlabel metal2 s 12810 12980 12918 13090 4 gnd
port 541 nsew
rlabel metal2 s 7818 5080 7926 5190 4 gnd
port 541 nsew
rlabel metal2 s 5802 10864 5910 10940 4 gnd
port 541 nsew
rlabel metal2 s 10794 9284 10902 9360 4 gnd
port 541 nsew
rlabel metal2 s 330 20660 438 20736 4 gnd
port 541 nsew
rlabel metal2 s 13290 13550 13398 13626 4 gnd
port 541 nsew
rlabel metal2 s 16554 1700 16662 1776 4 gnd
port 541 nsew
rlabel metal2 s 14058 13770 14166 13880 4 gnd
port 541 nsew
rlabel metal2 s 5322 15920 5430 15996 4 gnd
port 541 nsew
rlabel metal2 s 16554 14814 16662 14890 4 gnd
port 541 nsew
rlabel metal2 s 810 5870 918 5980 4 gnd
port 541 nsew
rlabel metal2 s 20778 13770 20886 13880 4 gnd
port 541 nsew
rlabel metal2 s 12042 9284 12150 9360 4 gnd
port 541 nsew
rlabel metal2 s 7818 2710 7926 2820 4 gnd
port 541 nsew
rlabel metal2 s 13290 9284 13398 9360 4 gnd
port 541 nsew
rlabel metal2 s 8298 1130 8406 1240 4 gnd
port 541 nsew
rlabel metal2 s 15306 8494 15414 8570 4 gnd
port 541 nsew
rlabel metal2 s 4554 1130 4662 1240 4 gnd
port 541 nsew
rlabel metal2 s 20778 21670 20886 21780 4 gnd
port 541 nsew
rlabel metal2 s 1578 21670 1686 21780 4 gnd
port 541 nsew
rlabel metal2 s 17802 23250 17910 23360 4 gnd
port 541 nsew
rlabel metal2 s 20778 19300 20886 19410 4 gnd
port 541 nsew
rlabel metal2 s 15306 24040 15414 24150 4 gnd
port 541 nsew
rlabel metal2 s 17034 20880 17142 20990 4 gnd
port 541 nsew
rlabel metal2 s 10794 2174 10902 2250 4 gnd
port 541 nsew
rlabel metal2 s 9066 18510 9174 18620 4 gnd
port 541 nsew
rlabel metal2 s 15786 3754 15894 3830 4 gnd
port 541 nsew
rlabel metal2 s 9546 13234 9654 13310 4 gnd
port 541 nsew
rlabel metal2 s 1578 11654 1686 11730 4 gnd
port 541 nsew
rlabel metal2 s 18282 8240 18390 8350 4 gnd
port 541 nsew
rlabel metal2 s 18282 2964 18390 3040 4 gnd
port 541 nsew
rlabel metal2 s 9546 17974 9654 18050 4 gnd
port 541 nsew
rlabel metal2 s 7818 8494 7926 8570 4 gnd
port 541 nsew
rlabel metal2 s 14058 11400 14166 11510 4 gnd
port 541 nsew
rlabel metal2 s 5322 10610 5430 10720 4 gnd
port 541 nsew
rlabel metal2 s 17034 5870 17142 5980 4 gnd
port 541 nsew
rlabel metal2 s 330 23250 438 23360 4 gnd
port 541 nsew
rlabel metal2 s 3306 21924 3414 22000 4 gnd
port 541 nsew
rlabel metal2 s 18282 18510 18390 18620 4 gnd
port 541 nsew
rlabel metal2 s 14538 25620 14646 25730 4 gnd
port 541 nsew
rlabel metal2 s 16554 5870 16662 5980 4 gnd
port 541 nsew
rlabel metal2 s 17802 2174 17910 2250 4 gnd
port 541 nsew
rlabel metal2 s 6570 5080 6678 5190 4 gnd
port 541 nsew
rlabel metal2 s 7818 17720 7926 17830 4 gnd
port 541 nsew
rlabel metal2 s 12042 12444 12150 12520 4 gnd
port 541 nsew
rlabel metal2 s 5322 25874 5430 25950 4 gnd
port 541 nsew
rlabel metal2 s 5322 20660 5430 20736 4 gnd
port 541 nsew
rlabel metal2 s 2826 120 2934 196 4 gnd
port 541 nsew
rlabel metal2 s 14538 910 14646 986 4 gnd
port 541 nsew
rlabel metal2 s 10794 1130 10902 1240 4 gnd
port 541 nsew
rlabel metal2 s 16554 10390 16662 10466 4 gnd
port 541 nsew
rlabel metal2 s 5322 20880 5430 20990 4 gnd
port 541 nsew
rlabel metal2 s 810 15604 918 15680 4 gnd
port 541 nsew
rlabel metal2 s 5802 10390 5910 10466 4 gnd
port 541 nsew
rlabel metal2 s 11562 4860 11670 4936 4 gnd
port 541 nsew
rlabel metal2 s 10794 910 10902 986 4 gnd
port 541 nsew
rlabel metal2 s 330 10610 438 10720 4 gnd
port 541 nsew
rlabel metal2 s 2826 22714 2934 22790 4 gnd
port 541 nsew
rlabel metal2 s 9546 2174 9654 2250 4 gnd
port 541 nsew
rlabel metal2 s 3306 7450 3414 7560 4 gnd
port 541 nsew
rlabel metal2 s 810 23820 918 23896 4 gnd
port 541 nsew
rlabel metal2 s 3306 22714 3414 22790 4 gnd
port 541 nsew
rlabel metal2 s 20778 9820 20886 9930 4 gnd
port 541 nsew
rlabel metal2 s 4074 5650 4182 5726 4 gnd
port 541 nsew
rlabel metal2 s 4074 594 4182 670 4 gnd
port 541 nsew
rlabel metal2 s 19530 25620 19638 25730 4 gnd
port 541 nsew
rlabel metal2 s 7050 25620 7158 25730 4 gnd
port 541 nsew
rlabel metal2 s 8298 1700 8406 1776 4 gnd
port 541 nsew
rlabel metal2 s 4074 16140 4182 16250 4 gnd
port 541 nsew
rlabel metal2 s 5322 120 5430 196 4 gnd
port 541 nsew
rlabel metal2 s 9546 340 9654 450 4 gnd
port 541 nsew
rlabel metal2 s 3306 340 3414 450 4 gnd
port 541 nsew
rlabel metal2 s 16554 16140 16662 16250 4 gnd
port 541 nsew
rlabel metal2 s 18282 11180 18390 11256 4 gnd
port 541 nsew
rlabel metal2 s 3306 12190 3414 12300 4 gnd
port 541 nsew
rlabel metal2 s 20778 17974 20886 18050 4 gnd
port 541 nsew
rlabel metal2 s 17802 9030 17910 9140 4 gnd
port 541 nsew
rlabel metal2 s 18282 17720 18390 17830 4 gnd
port 541 nsew
rlabel metal2 s 1578 1700 1686 1776 4 gnd
port 541 nsew
rlabel metal2 s 15786 20660 15894 20736 4 gnd
port 541 nsew
rlabel metal2 s 17802 15920 17910 15996 4 gnd
port 541 nsew
rlabel metal2 s 20778 7230 20886 7306 4 gnd
port 541 nsew
rlabel metal2 s 17802 8240 17910 8350 4 gnd
port 541 nsew
rlabel metal2 s 2058 20660 2166 20736 4 gnd
port 541 nsew
rlabel metal2 s 7818 23030 7926 23106 4 gnd
port 541 nsew
rlabel metal2 s 4074 24610 4182 24686 4 gnd
port 541 nsew
rlabel metal2 s 7818 17184 7926 17260 4 gnd
port 541 nsew
rlabel metal2 s 9546 23820 9654 23896 4 gnd
port 541 nsew
rlabel metal2 s 18282 16710 18390 16786 4 gnd
port 541 nsew
rlabel metal2 s 14058 4070 14166 4146 4 gnd
port 541 nsew
rlabel metal2 s 12810 1700 12918 1776 4 gnd
port 541 nsew
rlabel metal2 s 6570 10864 6678 10940 4 gnd
port 541 nsew
rlabel metal2 s 6570 19554 6678 19630 4 gnd
port 541 nsew
rlabel metal2 s 9066 17974 9174 18050 4 gnd
port 541 nsew
rlabel metal2 s 12042 21924 12150 22000 4 gnd
port 541 nsew
rlabel metal2 s 19050 13550 19158 13626 4 gnd
port 541 nsew
rlabel metal2 s 15306 4290 15414 4400 4 gnd
port 541 nsew
rlabel metal2 s 4074 8240 4182 8350 4 gnd
port 541 nsew
rlabel metal2 s 15786 25400 15894 25476 4 gnd
port 541 nsew
rlabel metal2 s 8298 14024 8406 14100 4 gnd
port 541 nsew
rlabel metal2 s 330 2490 438 2566 4 gnd
port 541 nsew
rlabel metal2 s 5802 5650 5910 5726 4 gnd
port 541 nsew
rlabel metal2 s 7818 8020 7926 8096 4 gnd
port 541 nsew
rlabel metal2 s 19050 24040 19158 24150 4 gnd
port 541 nsew
rlabel metal2 s 9546 24830 9654 24940 4 gnd
port 541 nsew
rlabel metal2 s 10314 4860 10422 4936 4 gnd
port 541 nsew
rlabel metal2 s 15786 10864 15894 10940 4 gnd
port 541 nsew
rlabel metal2 s 15306 23504 15414 23580 4 gnd
port 541 nsew
rlabel metal2 s 9066 18290 9174 18366 4 gnd
port 541 nsew
rlabel metal2 s 9066 23250 9174 23360 4 gnd
port 541 nsew
rlabel metal2 s 15786 20090 15894 20200 4 gnd
port 541 nsew
rlabel metal2 s 15306 13770 15414 13880 4 gnd
port 541 nsew
rlabel metal2 s 12042 5650 12150 5726 4 gnd
port 541 nsew
rlabel metal2 s 17034 17500 17142 17576 4 gnd
port 541 nsew
rlabel metal2 s 2058 15604 2166 15680 4 gnd
port 541 nsew
rlabel metal2 s 12810 340 12918 450 4 gnd
port 541 nsew
rlabel metal2 s 13290 24040 13398 24150 4 gnd
port 541 nsew
rlabel metal2 s 10794 6914 10902 6990 4 gnd
port 541 nsew
rlabel metal2 s 13290 15130 13398 15206 4 gnd
port 541 nsew
rlabel metal2 s 13290 13770 13398 13880 4 gnd
port 541 nsew
rlabel metal2 s 9546 17720 9654 17830 4 gnd
port 541 nsew
rlabel metal2 s 11562 8020 11670 8096 4 gnd
port 541 nsew
rlabel metal2 s 15306 9284 15414 9360 4 gnd
port 541 nsew
rlabel metal2 s 19050 2964 19158 3040 4 gnd
port 541 nsew
rlabel metal2 s 14058 20090 14166 20200 4 gnd
port 541 nsew
rlabel metal2 s 14538 12444 14646 12520 4 gnd
port 541 nsew
rlabel metal2 s 4554 9600 4662 9676 4 gnd
port 541 nsew
rlabel metal2 s 12810 2174 12918 2250 4 gnd
port 541 nsew
rlabel metal2 s 20778 24294 20886 24370 4 gnd
port 541 nsew
rlabel metal2 s 5322 19300 5430 19410 4 gnd
port 541 nsew
rlabel metal2 s 4554 18510 4662 18620 4 gnd
port 541 nsew
rlabel metal2 s 11562 11180 11670 11256 4 gnd
port 541 nsew
rlabel metal2 s 12042 6124 12150 6200 4 gnd
port 541 nsew
rlabel metal2 s 13290 120 13398 196 4 gnd
port 541 nsew
rlabel metal2 s 15306 6914 15414 6990 4 gnd
port 541 nsew
rlabel metal2 s 4074 11180 4182 11256 4 gnd
port 541 nsew
rlabel metal2 s 16554 14340 16662 14416 4 gnd
port 541 nsew
rlabel metal2 s 12042 20880 12150 20990 4 gnd
port 541 nsew
rlabel metal2 s 20298 4860 20406 4936 4 gnd
port 541 nsew
rlabel metal2 s 17034 19300 17142 19410 4 gnd
port 541 nsew
rlabel metal2 s 9066 23504 9174 23580 4 gnd
port 541 nsew
rlabel metal2 s 4554 20880 4662 20990 4 gnd
port 541 nsew
rlabel metal2 s 330 6124 438 6200 4 gnd
port 541 nsew
rlabel metal2 s 5322 3500 5430 3610 4 gnd
port 541 nsew
rlabel metal2 s 9066 2710 9174 2820 4 gnd
port 541 nsew
rlabel metal2 s 15786 19870 15894 19946 4 gnd
port 541 nsew
rlabel metal2 s 15786 19300 15894 19410 4 gnd
port 541 nsew
rlabel metal2 s 19050 6124 19158 6200 4 gnd
port 541 nsew
rlabel metal2 s 12810 14814 12918 14890 4 gnd
port 541 nsew
rlabel metal2 s 12042 22240 12150 22316 4 gnd
port 541 nsew
rlabel metal2 s 1578 12980 1686 13090 4 gnd
port 541 nsew
rlabel metal2 s 14058 2964 14166 3040 4 gnd
port 541 nsew
rlabel metal2 s 16554 13550 16662 13626 4 gnd
port 541 nsew
rlabel metal2 s 17034 13234 17142 13310 4 gnd
port 541 nsew
rlabel metal2 s 13290 14024 13398 14100 4 gnd
port 541 nsew
rlabel metal2 s 9546 14560 9654 14670 4 gnd
port 541 nsew
rlabel metal2 s 13290 7450 13398 7560 4 gnd
port 541 nsew
rlabel metal2 s 5322 4290 5430 4400 4 gnd
port 541 nsew
rlabel metal2 s 10314 19080 10422 19156 4 gnd
port 541 nsew
rlabel metal2 s 15306 22240 15414 22316 4 gnd
port 541 nsew
rlabel metal2 s 8298 12760 8406 12836 4 gnd
port 541 nsew
rlabel metal2 s 1578 5334 1686 5410 4 gnd
port 541 nsew
rlabel metal2 s 14538 9284 14646 9360 4 gnd
port 541 nsew
rlabel metal2 s 15306 7230 15414 7306 4 gnd
port 541 nsew
rlabel metal2 s 4554 19300 4662 19410 4 gnd
port 541 nsew
rlabel metal2 s 7050 7230 7158 7306 4 gnd
port 541 nsew
rlabel metal2 s 7050 4070 7158 4146 4 gnd
port 541 nsew
rlabel metal2 s 7050 2490 7158 2566 4 gnd
port 541 nsew
rlabel metal2 s 1578 25620 1686 25730 4 gnd
port 541 nsew
rlabel metal2 s 16554 25620 16662 25730 4 gnd
port 541 nsew
rlabel metal2 s 5802 15920 5910 15996 4 gnd
port 541 nsew
rlabel metal2 s 19530 24830 19638 24940 4 gnd
port 541 nsew
rlabel metal2 s 4554 15920 4662 15996 4 gnd
port 541 nsew
rlabel metal2 s 10314 23030 10422 23106 4 gnd
port 541 nsew
rlabel metal2 s 7050 21134 7158 21210 4 gnd
port 541 nsew
rlabel metal2 s 12042 23030 12150 23106 4 gnd
port 541 nsew
rlabel metal2 s 4554 16140 4662 16250 4 gnd
port 541 nsew
rlabel metal2 s 16554 10074 16662 10150 4 gnd
port 541 nsew
rlabel metal2 s 19050 19554 19158 19630 4 gnd
port 541 nsew
rlabel metal2 s 9546 21670 9654 21780 4 gnd
port 541 nsew
rlabel metal2 s 9546 910 9654 986 4 gnd
port 541 nsew
rlabel metal2 s 12042 6440 12150 6516 4 gnd
port 541 nsew
rlabel metal2 s 2058 9600 2166 9676 4 gnd
port 541 nsew
rlabel metal2 s 14538 20090 14646 20200 4 gnd
port 541 nsew
rlabel metal2 s 1578 910 1686 986 4 gnd
port 541 nsew
rlabel metal2 s 15306 13550 15414 13626 4 gnd
port 541 nsew
rlabel metal2 s 1578 15130 1686 15206 4 gnd
port 541 nsew
rlabel metal2 s 4554 13234 4662 13310 4 gnd
port 541 nsew
rlabel metal2 s 7818 10864 7926 10940 4 gnd
port 541 nsew
rlabel metal2 s 5322 13234 5430 13310 4 gnd
port 541 nsew
rlabel metal2 s 18282 11400 18390 11510 4 gnd
port 541 nsew
rlabel metal2 s 9546 5334 9654 5410 4 gnd
port 541 nsew
rlabel metal2 s 7818 594 7926 670 4 gnd
port 541 nsew
rlabel metal2 s 7050 4290 7158 4400 4 gnd
port 541 nsew
rlabel metal2 s 11562 7230 11670 7306 4 gnd
port 541 nsew
rlabel metal2 s 18282 22240 18390 22316 4 gnd
port 541 nsew
rlabel metal2 s 10794 21134 10902 21210 4 gnd
port 541 nsew
rlabel metal2 s 4554 13770 4662 13880 4 gnd
port 541 nsew
rlabel metal2 s 10794 17500 10902 17576 4 gnd
port 541 nsew
rlabel metal2 s 3306 19870 3414 19946 4 gnd
port 541 nsew
rlabel metal2 s 13290 21924 13398 22000 4 gnd
port 541 nsew
rlabel metal2 s 15306 22714 15414 22790 4 gnd
port 541 nsew
rlabel metal2 s 14058 23250 14166 23360 4 gnd
port 541 nsew
rlabel metal2 s 12810 21670 12918 21780 4 gnd
port 541 nsew
rlabel metal2 s 20778 4544 20886 4620 4 gnd
port 541 nsew
rlabel metal2 s 11562 12190 11670 12300 4 gnd
port 541 nsew
rlabel metal2 s 14058 10074 14166 10150 4 gnd
port 541 nsew
rlabel metal2 s 16554 11654 16662 11730 4 gnd
port 541 nsew
rlabel metal2 s 19530 1384 19638 1460 4 gnd
port 541 nsew
rlabel metal2 s 19050 7230 19158 7306 4 gnd
port 541 nsew
rlabel metal2 s 330 11970 438 12046 4 gnd
port 541 nsew
rlabel metal2 s 12042 22714 12150 22790 4 gnd
port 541 nsew
rlabel metal2 s 13290 5334 13398 5410 4 gnd
port 541 nsew
rlabel metal2 s 4554 19080 4662 19156 4 gnd
port 541 nsew
rlabel metal2 s 9066 14560 9174 14670 4 gnd
port 541 nsew
rlabel metal2 s 14538 6124 14646 6200 4 gnd
port 541 nsew
rlabel metal2 s 4074 25400 4182 25476 4 gnd
port 541 nsew
rlabel metal2 s 9546 14024 9654 14100 4 gnd
port 541 nsew
rlabel metal2 s 20298 9600 20406 9676 4 gnd
port 541 nsew
rlabel metal2 s 17034 24610 17142 24686 4 gnd
port 541 nsew
rlabel metal2 s 12810 19300 12918 19410 4 gnd
port 541 nsew
rlabel metal2 s 15306 4544 15414 4620 4 gnd
port 541 nsew
rlabel metal2 s 5322 23820 5430 23896 4 gnd
port 541 nsew
rlabel metal2 s 18282 24294 18390 24370 4 gnd
port 541 nsew
rlabel metal2 s 10794 9030 10902 9140 4 gnd
port 541 nsew
rlabel metal2 s 10794 17974 10902 18050 4 gnd
port 541 nsew
rlabel metal2 s 4554 20344 4662 20420 4 gnd
port 541 nsew
rlabel metal2 s 8298 21450 8406 21526 4 gnd
port 541 nsew
rlabel metal2 s 9546 20090 9654 20200 4 gnd
port 541 nsew
rlabel metal2 s 17034 17184 17142 17260 4 gnd
port 541 nsew
rlabel metal2 s 8298 11654 8406 11730 4 gnd
port 541 nsew
rlabel metal2 s 13290 594 13398 670 4 gnd
port 541 nsew
rlabel metal2 s 12042 2964 12150 3040 4 gnd
port 541 nsew
rlabel metal2 s 19050 11180 19158 11256 4 gnd
port 541 nsew
rlabel metal2 s 19050 7450 19158 7560 4 gnd
port 541 nsew
rlabel metal2 s 20298 910 20406 986 4 gnd
port 541 nsew
rlabel metal2 s 6570 17184 6678 17260 4 gnd
port 541 nsew
rlabel metal2 s 15306 16140 15414 16250 4 gnd
port 541 nsew
rlabel metal2 s 14058 16930 14166 17040 4 gnd
port 541 nsew
rlabel metal2 s 14058 910 14166 986 4 gnd
port 541 nsew
rlabel metal2 s 15306 25400 15414 25476 4 gnd
port 541 nsew
rlabel metal2 s 2058 21924 2166 22000 4 gnd
port 541 nsew
rlabel metal2 s 11562 25400 11670 25476 4 gnd
port 541 nsew
rlabel metal2 s 18282 1130 18390 1240 4 gnd
port 541 nsew
rlabel metal2 s 16554 24294 16662 24370 4 gnd
port 541 nsew
rlabel metal2 s 1578 6440 1686 6516 4 gnd
port 541 nsew
rlabel metal2 s 12810 22714 12918 22790 4 gnd
port 541 nsew
rlabel metal2 s 11562 9030 11670 9140 4 gnd
port 541 nsew
rlabel metal2 s 5322 15350 5430 15460 4 gnd
port 541 nsew
rlabel metal2 s 14538 18764 14646 18840 4 gnd
port 541 nsew
rlabel metal2 s 9546 16140 9654 16250 4 gnd
port 541 nsew
rlabel metal2 s 810 23250 918 23360 4 gnd
port 541 nsew
rlabel metal2 s 14538 2490 14646 2566 4 gnd
port 541 nsew
rlabel metal2 s 2826 21450 2934 21526 4 gnd
port 541 nsew
rlabel metal2 s 5802 24830 5910 24940 4 gnd
port 541 nsew
rlabel metal2 s 2826 22460 2934 22570 4 gnd
port 541 nsew
rlabel metal2 s 15786 8494 15894 8570 4 gnd
port 541 nsew
rlabel metal2 s 12810 2964 12918 3040 4 gnd
port 541 nsew
rlabel metal2 s 12042 17974 12150 18050 4 gnd
port 541 nsew
rlabel metal2 s 14058 22240 14166 22316 4 gnd
port 541 nsew
rlabel metal2 s 12810 8240 12918 8350 4 gnd
port 541 nsew
rlabel metal2 s 5322 5650 5430 5726 4 gnd
port 541 nsew
rlabel metal2 s 18282 14560 18390 14670 4 gnd
port 541 nsew
rlabel metal2 s 3306 4544 3414 4620 4 gnd
port 541 nsew
rlabel metal2 s 2058 8240 2166 8350 4 gnd
port 541 nsew
rlabel metal2 s 19050 8240 19158 8350 4 gnd
port 541 nsew
rlabel metal2 s 5802 12444 5910 12520 4 gnd
port 541 nsew
rlabel metal2 s 20298 11970 20406 12046 4 gnd
port 541 nsew
rlabel metal2 s 2826 3754 2934 3830 4 gnd
port 541 nsew
rlabel metal2 s 4554 16930 4662 17040 4 gnd
port 541 nsew
rlabel metal2 s 12810 594 12918 670 4 gnd
port 541 nsew
rlabel metal2 s 20298 14814 20406 14890 4 gnd
port 541 nsew
rlabel metal2 s 3306 18510 3414 18620 4 gnd
port 541 nsew
rlabel metal2 s 5802 19300 5910 19410 4 gnd
port 541 nsew
rlabel metal2 s 5802 8240 5910 8350 4 gnd
port 541 nsew
rlabel metal2 s 10794 10864 10902 10940 4 gnd
port 541 nsew
rlabel metal2 s 15306 7704 15414 7780 4 gnd
port 541 nsew
rlabel metal2 s 2826 12980 2934 13090 4 gnd
port 541 nsew
rlabel metal2 s 20778 11654 20886 11730 4 gnd
port 541 nsew
rlabel metal2 s 14058 5650 14166 5726 4 gnd
port 541 nsew
rlabel metal2 s 10794 19870 10902 19946 4 gnd
port 541 nsew
rlabel metal2 s 6570 15920 6678 15996 4 gnd
port 541 nsew
rlabel metal2 s 10314 1130 10422 1240 4 gnd
port 541 nsew
rlabel metal2 s 4554 22714 4662 22790 4 gnd
port 541 nsew
rlabel metal2 s 3306 8494 3414 8570 4 gnd
port 541 nsew
rlabel metal2 s 810 25084 918 25160 4 gnd
port 541 nsew
rlabel metal2 s 3306 25084 3414 25160 4 gnd
port 541 nsew
rlabel metal2 s 4074 1384 4182 1460 4 gnd
port 541 nsew
rlabel metal2 s 4554 24610 4662 24686 4 gnd
port 541 nsew
rlabel metal2 s 15306 2710 15414 2820 4 gnd
port 541 nsew
rlabel metal2 s 8298 19080 8406 19156 4 gnd
port 541 nsew
rlabel metal2 s 19050 5334 19158 5410 4 gnd
port 541 nsew
rlabel metal2 s 810 11654 918 11730 4 gnd
port 541 nsew
rlabel metal2 s 7818 21450 7926 21526 4 gnd
port 541 nsew
rlabel metal2 s 330 22240 438 22316 4 gnd
port 541 nsew
rlabel metal2 s 19530 6660 19638 6770 4 gnd
port 541 nsew
rlabel metal2 s 10794 23820 10902 23896 4 gnd
port 541 nsew
rlabel metal2 s 20778 20344 20886 20420 4 gnd
port 541 nsew
rlabel metal2 s 6570 5650 6678 5726 4 gnd
port 541 nsew
rlabel metal2 s 5802 4544 5910 4620 4 gnd
port 541 nsew
rlabel metal2 s 6570 2710 6678 2820 4 gnd
port 541 nsew
rlabel metal2 s 4074 13550 4182 13626 4 gnd
port 541 nsew
rlabel metal2 s 9066 1700 9174 1776 4 gnd
port 541 nsew
rlabel metal2 s 9546 7704 9654 7780 4 gnd
port 541 nsew
rlabel metal2 s 5322 10864 5430 10940 4 gnd
port 541 nsew
rlabel metal2 s 330 23504 438 23580 4 gnd
port 541 nsew
rlabel metal2 s 2058 24830 2166 24940 4 gnd
port 541 nsew
rlabel metal2 s 330 5870 438 5980 4 gnd
port 541 nsew
rlabel metal2 s 2826 11180 2934 11256 4 gnd
port 541 nsew
rlabel metal2 s 10794 3754 10902 3830 4 gnd
port 541 nsew
rlabel metal2 s 14538 5334 14646 5410 4 gnd
port 541 nsew
rlabel metal2 s 5802 20660 5910 20736 4 gnd
port 541 nsew
rlabel metal2 s 5322 16710 5430 16786 4 gnd
port 541 nsew
rlabel metal2 s 4074 7704 4182 7780 4 gnd
port 541 nsew
rlabel metal2 s 12810 120 12918 196 4 gnd
port 541 nsew
rlabel metal2 s 6570 23820 6678 23896 4 gnd
port 541 nsew
rlabel metal2 s 16554 16930 16662 17040 4 gnd
port 541 nsew
rlabel metal2 s 7818 21670 7926 21780 4 gnd
port 541 nsew
rlabel metal2 s 16554 12760 16662 12836 4 gnd
port 541 nsew
rlabel metal2 s 20778 9284 20886 9360 4 gnd
port 541 nsew
rlabel metal2 s 5322 24830 5430 24940 4 gnd
port 541 nsew
rlabel metal2 s 12042 12190 12150 12300 4 gnd
port 541 nsew
rlabel metal2 s 8298 9030 8406 9140 4 gnd
port 541 nsew
rlabel metal2 s 11562 25620 11670 25730 4 gnd
port 541 nsew
rlabel metal2 s 2058 21670 2166 21780 4 gnd
port 541 nsew
rlabel metal2 s 6570 11400 6678 11510 4 gnd
port 541 nsew
rlabel metal2 s 20298 20090 20406 20200 4 gnd
port 541 nsew
rlabel metal2 s 6570 15604 6678 15680 4 gnd
port 541 nsew
rlabel metal2 s 5802 17184 5910 17260 4 gnd
port 541 nsew
rlabel metal2 s 12042 3500 12150 3610 4 gnd
port 541 nsew
rlabel metal2 s 15306 18764 15414 18840 4 gnd
port 541 nsew
rlabel metal2 s 1578 10074 1686 10150 4 gnd
port 541 nsew
rlabel metal2 s 3306 15130 3414 15206 4 gnd
port 541 nsew
rlabel metal2 s 7050 21924 7158 22000 4 gnd
port 541 nsew
rlabel metal2 s 810 2710 918 2820 4 gnd
port 541 nsew
rlabel metal2 s 17034 120 17142 196 4 gnd
port 541 nsew
rlabel metal2 s 8298 24830 8406 24940 4 gnd
port 541 nsew
rlabel metal2 s 9066 6440 9174 6516 4 gnd
port 541 nsew
rlabel metal2 s 9066 7450 9174 7560 4 gnd
port 541 nsew
rlabel metal2 s 1578 6914 1686 6990 4 gnd
port 541 nsew
rlabel metal2 s 2058 4860 2166 4936 4 gnd
port 541 nsew
rlabel metal2 s 9066 10610 9174 10720 4 gnd
port 541 nsew
rlabel metal2 s 12810 25620 12918 25730 4 gnd
port 541 nsew
rlabel metal2 s 20778 21134 20886 21210 4 gnd
port 541 nsew
rlabel metal2 s 6570 8020 6678 8096 4 gnd
port 541 nsew
rlabel metal2 s 20778 10074 20886 10150 4 gnd
port 541 nsew
rlabel metal2 s 18282 16930 18390 17040 4 gnd
port 541 nsew
rlabel metal2 s 14538 9030 14646 9140 4 gnd
port 541 nsew
rlabel metal2 s 15786 11654 15894 11730 4 gnd
port 541 nsew
rlabel metal2 s 10794 20090 10902 20200 4 gnd
port 541 nsew
rlabel metal2 s 330 1920 438 2030 4 gnd
port 541 nsew
rlabel metal2 s 17802 2710 17910 2820 4 gnd
port 541 nsew
rlabel metal2 s 9546 4860 9654 4936 4 gnd
port 541 nsew
rlabel metal2 s 20778 22240 20886 22316 4 gnd
port 541 nsew
rlabel metal2 s 15306 12190 15414 12300 4 gnd
port 541 nsew
rlabel metal2 s 8298 5080 8406 5190 4 gnd
port 541 nsew
rlabel metal2 s 4554 8240 4662 8350 4 gnd
port 541 nsew
rlabel metal2 s 20298 6660 20406 6770 4 gnd
port 541 nsew
rlabel metal2 s 9546 11654 9654 11730 4 gnd
port 541 nsew
rlabel metal2 s 3306 13550 3414 13626 4 gnd
port 541 nsew
rlabel metal2 s 12810 23030 12918 23106 4 gnd
port 541 nsew
rlabel metal2 s 330 25084 438 25160 4 gnd
port 541 nsew
rlabel metal2 s 19050 21670 19158 21780 4 gnd
port 541 nsew
rlabel metal2 s 11562 20880 11670 20990 4 gnd
port 541 nsew
rlabel metal2 s 20298 22714 20406 22790 4 gnd
port 541 nsew
rlabel metal2 s 20778 14814 20886 14890 4 gnd
port 541 nsew
rlabel metal2 s 11562 19300 11670 19410 4 gnd
port 541 nsew
rlabel metal2 s 5322 10074 5430 10150 4 gnd
port 541 nsew
rlabel metal2 s 14538 17184 14646 17260 4 gnd
port 541 nsew
rlabel metal2 s 810 2964 918 3040 4 gnd
port 541 nsew
rlabel metal2 s 12042 6660 12150 6770 4 gnd
port 541 nsew
rlabel metal2 s 4554 3500 4662 3610 4 gnd
port 541 nsew
rlabel metal2 s 6570 15130 6678 15206 4 gnd
port 541 nsew
rlabel metal2 s 10314 21134 10422 21210 4 gnd
port 541 nsew
rlabel metal2 s 5802 7230 5910 7306 4 gnd
port 541 nsew
rlabel metal2 s 9546 4070 9654 4146 4 gnd
port 541 nsew
rlabel metal2 s 810 18510 918 18620 4 gnd
port 541 nsew
rlabel metal2 s 17034 6914 17142 6990 4 gnd
port 541 nsew
rlabel metal2 s 12042 8240 12150 8350 4 gnd
port 541 nsew
rlabel metal2 s 19530 18764 19638 18840 4 gnd
port 541 nsew
rlabel metal2 s 14538 25084 14646 25160 4 gnd
port 541 nsew
rlabel metal2 s 12042 12980 12150 13090 4 gnd
port 541 nsew
rlabel metal2 s 11562 15604 11670 15680 4 gnd
port 541 nsew
rlabel metal2 s 4554 340 4662 450 4 gnd
port 541 nsew
rlabel metal2 s 5322 24610 5430 24686 4 gnd
port 541 nsew
rlabel metal2 s 7050 10610 7158 10720 4 gnd
port 541 nsew
rlabel metal2 s 19050 16140 19158 16250 4 gnd
port 541 nsew
rlabel metal2 s 6570 9030 6678 9140 4 gnd
port 541 nsew
rlabel metal2 s 18282 7450 18390 7560 4 gnd
port 541 nsew
rlabel metal2 s 10794 15350 10902 15460 4 gnd
port 541 nsew
rlabel metal2 s 9066 15130 9174 15206 4 gnd
port 541 nsew
rlabel metal2 s 15306 22460 15414 22570 4 gnd
port 541 nsew
rlabel metal2 s 17802 13234 17910 13310 4 gnd
port 541 nsew
rlabel metal2 s 19530 10864 19638 10940 4 gnd
port 541 nsew
rlabel metal2 s 5322 4860 5430 4936 4 gnd
port 541 nsew
rlabel metal2 s 9066 24830 9174 24940 4 gnd
port 541 nsew
rlabel metal2 s 4554 7450 4662 7560 4 gnd
port 541 nsew
rlabel metal2 s 18282 19870 18390 19946 4 gnd
port 541 nsew
rlabel metal2 s 5802 11400 5910 11510 4 gnd
port 541 nsew
rlabel metal2 s 17034 10610 17142 10720 4 gnd
port 541 nsew
rlabel metal2 s 20778 22714 20886 22790 4 gnd
port 541 nsew
rlabel metal2 s 20778 5080 20886 5190 4 gnd
port 541 nsew
rlabel metal2 s 19530 25874 19638 25950 4 gnd
port 541 nsew
rlabel metal2 s 5802 24040 5910 24150 4 gnd
port 541 nsew
rlabel metal2 s 10314 5870 10422 5980 4 gnd
port 541 nsew
rlabel metal2 s 9066 23030 9174 23106 4 gnd
port 541 nsew
rlabel metal2 s 10794 12980 10902 13090 4 gnd
port 541 nsew
rlabel metal2 s 1578 12444 1686 12520 4 gnd
port 541 nsew
rlabel metal2 s 4554 14024 4662 14100 4 gnd
port 541 nsew
rlabel metal2 s 7818 18510 7926 18620 4 gnd
port 541 nsew
rlabel metal2 s 5802 8810 5910 8886 4 gnd
port 541 nsew
rlabel metal2 s 7818 4544 7926 4620 4 gnd
port 541 nsew
rlabel metal2 s 14058 4860 14166 4936 4 gnd
port 541 nsew
rlabel metal2 s 6570 12190 6678 12300 4 gnd
port 541 nsew
rlabel metal2 s 20778 8810 20886 8886 4 gnd
port 541 nsew
rlabel metal2 s 12810 23820 12918 23896 4 gnd
port 541 nsew
rlabel metal2 s 810 17974 918 18050 4 gnd
port 541 nsew
rlabel metal2 s 2826 12444 2934 12520 4 gnd
port 541 nsew
rlabel metal2 s 7818 21924 7926 22000 4 gnd
port 541 nsew
rlabel metal2 s 7050 8810 7158 8886 4 gnd
port 541 nsew
rlabel metal2 s 3306 14024 3414 14100 4 gnd
port 541 nsew
rlabel metal2 s 11562 12760 11670 12836 4 gnd
port 541 nsew
rlabel metal2 s 1578 22714 1686 22790 4 gnd
port 541 nsew
rlabel metal2 s 18282 20880 18390 20990 4 gnd
port 541 nsew
rlabel metal2 s 20298 2490 20406 2566 4 gnd
port 541 nsew
rlabel metal2 s 10794 17720 10902 17830 4 gnd
port 541 nsew
rlabel metal2 s 10314 3280 10422 3356 4 gnd
port 541 nsew
rlabel metal2 s 17034 14814 17142 14890 4 gnd
port 541 nsew
rlabel metal2 s 19050 8810 19158 8886 4 gnd
port 541 nsew
rlabel metal2 s 18282 19554 18390 19630 4 gnd
port 541 nsew
rlabel metal2 s 5802 4070 5910 4146 4 gnd
port 541 nsew
rlabel metal2 s 14058 1130 14166 1240 4 gnd
port 541 nsew
rlabel metal2 s 7818 21134 7926 21210 4 gnd
port 541 nsew
rlabel metal2 s 20298 17184 20406 17260 4 gnd
port 541 nsew
rlabel metal2 s 330 10864 438 10940 4 gnd
port 541 nsew
rlabel metal2 s 8298 4070 8406 4146 4 gnd
port 541 nsew
rlabel metal2 s 14058 15604 14166 15680 4 gnd
port 541 nsew
rlabel metal2 s 14538 23250 14646 23360 4 gnd
port 541 nsew
rlabel metal2 s 330 19870 438 19946 4 gnd
port 541 nsew
rlabel metal2 s 19530 13234 19638 13310 4 gnd
port 541 nsew
rlabel metal2 s 13290 11654 13398 11730 4 gnd
port 541 nsew
rlabel metal2 s 12042 17720 12150 17830 4 gnd
port 541 nsew
rlabel metal2 s 6570 24610 6678 24686 4 gnd
port 541 nsew
rlabel metal2 s 810 24040 918 24150 4 gnd
port 541 nsew
rlabel metal2 s 2058 3500 2166 3610 4 gnd
port 541 nsew
rlabel metal2 s 6570 10390 6678 10466 4 gnd
port 541 nsew
rlabel metal2 s 5802 6124 5910 6200 4 gnd
port 541 nsew
rlabel metal2 s 19530 16140 19638 16250 4 gnd
port 541 nsew
rlabel metal2 s 17034 23820 17142 23896 4 gnd
port 541 nsew
rlabel metal2 s 9546 19554 9654 19630 4 gnd
port 541 nsew
rlabel metal2 s 20778 14024 20886 14100 4 gnd
port 541 nsew
rlabel metal2 s 9066 5870 9174 5980 4 gnd
port 541 nsew
rlabel metal2 s 15786 16930 15894 17040 4 gnd
port 541 nsew
rlabel metal2 s 14538 22714 14646 22790 4 gnd
port 541 nsew
rlabel metal2 s 2826 19870 2934 19946 4 gnd
port 541 nsew
rlabel metal2 s 3306 23030 3414 23106 4 gnd
port 541 nsew
rlabel metal2 s 15786 18290 15894 18366 4 gnd
port 541 nsew
rlabel metal2 s 14538 8240 14646 8350 4 gnd
port 541 nsew
rlabel metal2 s 15306 11180 15414 11256 4 gnd
port 541 nsew
rlabel metal2 s 9066 1920 9174 2030 4 gnd
port 541 nsew
rlabel metal2 s 810 9820 918 9930 4 gnd
port 541 nsew
rlabel metal2 s 10794 24294 10902 24370 4 gnd
port 541 nsew
rlabel metal2 s 19050 22240 19158 22316 4 gnd
port 541 nsew
rlabel metal2 s 2058 9284 2166 9360 4 gnd
port 541 nsew
rlabel metal2 s 12042 18510 12150 18620 4 gnd
port 541 nsew
rlabel metal2 s 15786 10610 15894 10720 4 gnd
port 541 nsew
rlabel metal2 s 7818 10390 7926 10466 4 gnd
port 541 nsew
rlabel metal2 s 2826 21670 2934 21780 4 gnd
port 541 nsew
rlabel metal2 s 15306 17974 15414 18050 4 gnd
port 541 nsew
rlabel metal2 s 18282 4544 18390 4620 4 gnd
port 541 nsew
rlabel metal2 s 7050 9030 7158 9140 4 gnd
port 541 nsew
rlabel metal2 s 18282 910 18390 986 4 gnd
port 541 nsew
rlabel metal2 s 330 18764 438 18840 4 gnd
port 541 nsew
rlabel metal2 s 20778 19554 20886 19630 4 gnd
port 541 nsew
rlabel metal2 s 2826 23250 2934 23360 4 gnd
port 541 nsew
rlabel metal2 s 7050 23030 7158 23106 4 gnd
port 541 nsew
rlabel metal2 s 8298 21670 8406 21780 4 gnd
port 541 nsew
rlabel metal2 s 6570 8494 6678 8570 4 gnd
port 541 nsew
rlabel metal2 s 2826 24830 2934 24940 4 gnd
port 541 nsew
rlabel metal2 s 8298 14340 8406 14416 4 gnd
port 541 nsew
rlabel metal2 s 14538 11400 14646 11510 4 gnd
port 541 nsew
rlabel metal2 s 19530 6440 19638 6516 4 gnd
port 541 nsew
rlabel metal2 s 330 18510 438 18620 4 gnd
port 541 nsew
rlabel metal2 s 17802 1130 17910 1240 4 gnd
port 541 nsew
rlabel metal2 s 10794 1920 10902 2030 4 gnd
port 541 nsew
rlabel metal2 s 20778 14340 20886 14416 4 gnd
port 541 nsew
rlabel metal2 s 3306 8810 3414 8886 4 gnd
port 541 nsew
rlabel metal2 s 12810 11180 12918 11256 4 gnd
port 541 nsew
rlabel metal2 s 4554 5650 4662 5726 4 gnd
port 541 nsew
rlabel metal2 s 9546 9030 9654 9140 4 gnd
port 541 nsew
rlabel metal2 s 10314 20344 10422 20420 4 gnd
port 541 nsew
rlabel metal2 s 3306 2174 3414 2250 4 gnd
port 541 nsew
rlabel metal2 s 810 17500 918 17576 4 gnd
port 541 nsew
rlabel metal2 s 10794 13550 10902 13626 4 gnd
port 541 nsew
rlabel metal2 s 17034 24294 17142 24370 4 gnd
port 541 nsew
rlabel metal2 s 11562 910 11670 986 4 gnd
port 541 nsew
rlabel metal2 s 7050 910 7158 986 4 gnd
port 541 nsew
rlabel metal2 s 4554 2174 4662 2250 4 gnd
port 541 nsew
rlabel metal2 s 4074 15130 4182 15206 4 gnd
port 541 nsew
rlabel metal2 s 5802 14340 5910 14416 4 gnd
port 541 nsew
rlabel metal2 s 9546 15130 9654 15206 4 gnd
port 541 nsew
rlabel metal2 s 15786 11970 15894 12046 4 gnd
port 541 nsew
rlabel metal2 s 810 22460 918 22570 4 gnd
port 541 nsew
rlabel metal2 s 4074 23250 4182 23360 4 gnd
port 541 nsew
rlabel metal2 s 11562 16394 11670 16470 4 gnd
port 541 nsew
rlabel metal2 s 6570 3500 6678 3610 4 gnd
port 541 nsew
rlabel metal2 s 19050 22460 19158 22570 4 gnd
port 541 nsew
rlabel metal2 s 12810 18510 12918 18620 4 gnd
port 541 nsew
rlabel metal2 s 9066 20660 9174 20736 4 gnd
port 541 nsew
rlabel metal2 s 2058 2964 2166 3040 4 gnd
port 541 nsew
rlabel metal2 s 11562 14560 11670 14670 4 gnd
port 541 nsew
rlabel metal2 s 10314 20660 10422 20736 4 gnd
port 541 nsew
rlabel metal2 s 20298 22240 20406 22316 4 gnd
port 541 nsew
rlabel metal2 s 5802 21450 5910 21526 4 gnd
port 541 nsew
rlabel metal2 s 4074 6440 4182 6516 4 gnd
port 541 nsew
rlabel metal2 s 2058 5334 2166 5410 4 gnd
port 541 nsew
rlabel metal2 s 20298 8810 20406 8886 4 gnd
port 541 nsew
rlabel metal2 s 10794 22460 10902 22570 4 gnd
port 541 nsew
rlabel metal2 s 15786 23250 15894 23360 4 gnd
port 541 nsew
rlabel metal2 s 9066 5334 9174 5410 4 gnd
port 541 nsew
rlabel metal2 s 15786 4070 15894 4146 4 gnd
port 541 nsew
rlabel metal2 s 3306 11180 3414 11256 4 gnd
port 541 nsew
rlabel metal2 s 10794 18510 10902 18620 4 gnd
port 541 nsew
rlabel metal2 s 19050 15130 19158 15206 4 gnd
port 541 nsew
rlabel metal2 s 3306 14814 3414 14890 4 gnd
port 541 nsew
rlabel metal2 s 9546 6440 9654 6516 4 gnd
port 541 nsew
rlabel metal2 s 12042 10610 12150 10720 4 gnd
port 541 nsew
rlabel metal2 s 15786 24830 15894 24940 4 gnd
port 541 nsew
rlabel metal2 s 11562 24294 11670 24370 4 gnd
port 541 nsew
rlabel metal2 s 15306 3754 15414 3830 4 gnd
port 541 nsew
rlabel metal2 s 8298 20880 8406 20990 4 gnd
port 541 nsew
rlabel metal2 s 1578 2964 1686 3040 4 gnd
port 541 nsew
rlabel metal2 s 8298 11400 8406 11510 4 gnd
port 541 nsew
rlabel metal2 s 17802 5334 17910 5410 4 gnd
port 541 nsew
rlabel metal2 s 2826 18510 2934 18620 4 gnd
port 541 nsew
rlabel metal2 s 19050 340 19158 450 4 gnd
port 541 nsew
rlabel metal2 s 330 15130 438 15206 4 gnd
port 541 nsew
rlabel metal2 s 12042 15920 12150 15996 4 gnd
port 541 nsew
rlabel metal2 s 17802 7704 17910 7780 4 gnd
port 541 nsew
rlabel metal2 s 15786 10074 15894 10150 4 gnd
port 541 nsew
rlabel metal2 s 10314 23820 10422 23896 4 gnd
port 541 nsew
rlabel metal2 s 7050 20344 7158 20420 4 gnd
port 541 nsew
rlabel metal2 s 16554 7230 16662 7306 4 gnd
port 541 nsew
rlabel metal2 s 5322 1130 5430 1240 4 gnd
port 541 nsew
rlabel metal2 s 1578 8020 1686 8096 4 gnd
port 541 nsew
rlabel metal2 s 9546 22714 9654 22790 4 gnd
port 541 nsew
rlabel metal2 s 19530 19870 19638 19946 4 gnd
port 541 nsew
rlabel metal2 s 5322 8020 5430 8096 4 gnd
port 541 nsew
rlabel metal2 s 15306 6124 15414 6200 4 gnd
port 541 nsew
rlabel metal2 s 20778 11400 20886 11510 4 gnd
port 541 nsew
rlabel metal2 s 10794 10074 10902 10150 4 gnd
port 541 nsew
rlabel metal2 s 9066 10074 9174 10150 4 gnd
port 541 nsew
rlabel metal2 s 11562 10074 11670 10150 4 gnd
port 541 nsew
rlabel metal2 s 15306 21670 15414 21780 4 gnd
port 541 nsew
rlabel metal2 s 14058 20880 14166 20990 4 gnd
port 541 nsew
rlabel metal2 s 16554 21134 16662 21210 4 gnd
port 541 nsew
rlabel metal2 s 11562 17720 11670 17830 4 gnd
port 541 nsew
rlabel metal2 s 13290 23030 13398 23106 4 gnd
port 541 nsew
rlabel metal2 s 4074 20660 4182 20736 4 gnd
port 541 nsew
rlabel metal2 s 19530 910 19638 986 4 gnd
port 541 nsew
rlabel metal2 s 19530 2174 19638 2250 4 gnd
port 541 nsew
rlabel metal2 s 9066 8810 9174 8886 4 gnd
port 541 nsew
rlabel metal2 s 1578 3754 1686 3830 4 gnd
port 541 nsew
rlabel metal2 s 1578 594 1686 670 4 gnd
port 541 nsew
rlabel metal2 s 9546 11970 9654 12046 4 gnd
port 541 nsew
rlabel metal2 s 2058 18290 2166 18366 4 gnd
port 541 nsew
rlabel metal2 s 9066 25620 9174 25730 4 gnd
port 541 nsew
rlabel metal2 s 14058 24610 14166 24686 4 gnd
port 541 nsew
rlabel metal2 s 1578 11400 1686 11510 4 gnd
port 541 nsew
rlabel metal2 s 4074 5334 4182 5410 4 gnd
port 541 nsew
rlabel metal2 s 4554 8810 4662 8886 4 gnd
port 541 nsew
rlabel metal2 s 1578 19080 1686 19156 4 gnd
port 541 nsew
rlabel metal2 s 8298 25084 8406 25160 4 gnd
port 541 nsew
rlabel metal2 s 9066 19080 9174 19156 4 gnd
port 541 nsew
rlabel metal2 s 17802 24610 17910 24686 4 gnd
port 541 nsew
rlabel metal2 s 2058 11180 2166 11256 4 gnd
port 541 nsew
rlabel metal2 s 15786 13550 15894 13626 4 gnd
port 541 nsew
rlabel metal2 s 2058 21134 2166 21210 4 gnd
port 541 nsew
rlabel metal2 s 20778 8020 20886 8096 4 gnd
port 541 nsew
rlabel metal2 s 15306 11654 15414 11730 4 gnd
port 541 nsew
rlabel metal2 s 13290 23504 13398 23580 4 gnd
port 541 nsew
rlabel metal2 s 15306 24830 15414 24940 4 gnd
port 541 nsew
rlabel metal2 s 330 340 438 450 4 gnd
port 541 nsew
rlabel metal2 s 3306 16140 3414 16250 4 gnd
port 541 nsew
rlabel metal2 s 5322 5080 5430 5190 4 gnd
port 541 nsew
rlabel metal2 s 15306 5334 15414 5410 4 gnd
port 541 nsew
rlabel metal2 s 5322 5870 5430 5980 4 gnd
port 541 nsew
rlabel metal2 s 19050 9030 19158 9140 4 gnd
port 541 nsew
rlabel metal2 s 15306 910 15414 986 4 gnd
port 541 nsew
rlabel metal2 s 5322 21450 5430 21526 4 gnd
port 541 nsew
rlabel metal2 s 5802 4290 5910 4400 4 gnd
port 541 nsew
rlabel metal2 s 12810 15920 12918 15996 4 gnd
port 541 nsew
rlabel metal2 s 6570 11970 6678 12046 4 gnd
port 541 nsew
rlabel metal2 s 14538 12190 14646 12300 4 gnd
port 541 nsew
rlabel metal2 s 17802 11400 17910 11510 4 gnd
port 541 nsew
rlabel metal2 s 16554 4544 16662 4620 4 gnd
port 541 nsew
rlabel metal2 s 7050 17720 7158 17830 4 gnd
port 541 nsew
rlabel metal2 s 11562 20660 11670 20736 4 gnd
port 541 nsew
rlabel metal2 s 9066 22460 9174 22570 4 gnd
port 541 nsew
rlabel metal2 s 2058 16930 2166 17040 4 gnd
port 541 nsew
rlabel metal2 s 12042 10864 12150 10940 4 gnd
port 541 nsew
rlabel metal2 s 4554 9820 4662 9930 4 gnd
port 541 nsew
rlabel metal2 s 6570 4290 6678 4400 4 gnd
port 541 nsew
rlabel metal2 s 12042 9600 12150 9676 4 gnd
port 541 nsew
rlabel metal2 s 12810 19870 12918 19946 4 gnd
port 541 nsew
rlabel metal2 s 11562 14024 11670 14100 4 gnd
port 541 nsew
rlabel metal2 s 5322 23030 5430 23106 4 gnd
port 541 nsew
rlabel metal2 s 15786 7450 15894 7560 4 gnd
port 541 nsew
rlabel metal2 s 8298 15604 8406 15680 4 gnd
port 541 nsew
rlabel metal2 s 4074 21450 4182 21526 4 gnd
port 541 nsew
rlabel metal2 s 4554 6440 4662 6516 4 gnd
port 541 nsew
rlabel metal2 s 12810 7450 12918 7560 4 gnd
port 541 nsew
rlabel metal2 s 5322 18764 5430 18840 4 gnd
port 541 nsew
rlabel metal2 s 10314 6914 10422 6990 4 gnd
port 541 nsew
rlabel metal2 s 16554 17500 16662 17576 4 gnd
port 541 nsew
rlabel metal2 s 20778 22460 20886 22570 4 gnd
port 541 nsew
rlabel metal2 s 12042 19080 12150 19156 4 gnd
port 541 nsew
rlabel metal2 s 3306 16930 3414 17040 4 gnd
port 541 nsew
rlabel metal2 s 13290 1920 13398 2030 4 gnd
port 541 nsew
rlabel metal2 s 14058 4544 14166 4620 4 gnd
port 541 nsew
rlabel metal2 s 4074 10074 4182 10150 4 gnd
port 541 nsew
rlabel metal2 s 4074 16710 4182 16786 4 gnd
port 541 nsew
rlabel metal2 s 20298 17974 20406 18050 4 gnd
port 541 nsew
rlabel metal2 s 7818 19870 7926 19946 4 gnd
port 541 nsew
rlabel metal2 s 13290 20660 13398 20736 4 gnd
port 541 nsew
rlabel metal2 s 10314 120 10422 196 4 gnd
port 541 nsew
rlabel metal2 s 3306 3500 3414 3610 4 gnd
port 541 nsew
rlabel metal2 s 7050 12760 7158 12836 4 gnd
port 541 nsew
rlabel metal2 s 7818 24294 7926 24370 4 gnd
port 541 nsew
rlabel metal2 s 1578 6660 1686 6770 4 gnd
port 541 nsew
rlabel metal2 s 18282 2710 18390 2820 4 gnd
port 541 nsew
rlabel metal2 s 13290 12980 13398 13090 4 gnd
port 541 nsew
rlabel metal2 s 330 20344 438 20420 4 gnd
port 541 nsew
rlabel metal2 s 11562 3280 11670 3356 4 gnd
port 541 nsew
rlabel metal2 s 9066 16140 9174 16250 4 gnd
port 541 nsew
rlabel metal2 s 19530 24040 19638 24150 4 gnd
port 541 nsew
rlabel metal2 s 810 25400 918 25476 4 gnd
port 541 nsew
rlabel metal2 s 2826 25874 2934 25950 4 gnd
port 541 nsew
rlabel metal2 s 18282 24610 18390 24686 4 gnd
port 541 nsew
rlabel metal2 s 12042 120 12150 196 4 gnd
port 541 nsew
rlabel metal2 s 17802 2964 17910 3040 4 gnd
port 541 nsew
rlabel metal2 s 14058 14340 14166 14416 4 gnd
port 541 nsew
rlabel metal2 s 12042 11970 12150 12046 4 gnd
port 541 nsew
rlabel metal2 s 20778 5870 20886 5980 4 gnd
port 541 nsew
rlabel metal2 s 4074 4290 4182 4400 4 gnd
port 541 nsew
rlabel metal2 s 12042 20090 12150 20200 4 gnd
port 541 nsew
rlabel metal2 s 11562 5080 11670 5190 4 gnd
port 541 nsew
rlabel metal2 s 2826 24610 2934 24686 4 gnd
port 541 nsew
rlabel metal2 s 18282 22460 18390 22570 4 gnd
port 541 nsew
rlabel metal2 s 12810 14340 12918 14416 4 gnd
port 541 nsew
rlabel metal2 s 4074 11970 4182 12046 4 gnd
port 541 nsew
rlabel metal2 s 14538 1130 14646 1240 4 gnd
port 541 nsew
rlabel metal2 s 20778 20880 20886 20990 4 gnd
port 541 nsew
rlabel metal2 s 4074 6660 4182 6770 4 gnd
port 541 nsew
rlabel metal2 s 10794 4290 10902 4400 4 gnd
port 541 nsew
rlabel metal2 s 7050 17184 7158 17260 4 gnd
port 541 nsew
rlabel metal2 s 20778 17500 20886 17576 4 gnd
port 541 nsew
rlabel metal2 s 7050 21450 7158 21526 4 gnd
port 541 nsew
rlabel metal2 s 6570 13234 6678 13310 4 gnd
port 541 nsew
rlabel metal2 s 4074 18764 4182 18840 4 gnd
port 541 nsew
rlabel metal2 s 2826 23504 2934 23580 4 gnd
port 541 nsew
rlabel metal2 s 5802 120 5910 196 4 gnd
port 541 nsew
rlabel metal2 s 8298 5870 8406 5980 4 gnd
port 541 nsew
rlabel metal2 s 10314 910 10422 986 4 gnd
port 541 nsew
rlabel metal2 s 13290 17720 13398 17830 4 gnd
port 541 nsew
rlabel metal2 s 10314 17720 10422 17830 4 gnd
port 541 nsew
rlabel metal2 s 1578 16710 1686 16786 4 gnd
port 541 nsew
rlabel metal2 s 14058 15350 14166 15460 4 gnd
port 541 nsew
rlabel metal2 s 4074 2174 4182 2250 4 gnd
port 541 nsew
rlabel metal2 s 10794 5080 10902 5190 4 gnd
port 541 nsew
rlabel metal2 s 14538 6660 14646 6770 4 gnd
port 541 nsew
rlabel metal2 s 810 12444 918 12520 4 gnd
port 541 nsew
rlabel metal2 s 15786 1130 15894 1240 4 gnd
port 541 nsew
rlabel metal2 s 6570 594 6678 670 4 gnd
port 541 nsew
rlabel metal2 s 7818 20090 7926 20200 4 gnd
port 541 nsew
rlabel metal2 s 14058 3754 14166 3830 4 gnd
port 541 nsew
rlabel metal2 s 15306 20090 15414 20200 4 gnd
port 541 nsew
rlabel metal2 s 9546 11400 9654 11510 4 gnd
port 541 nsew
rlabel metal2 s 16554 20344 16662 20420 4 gnd
port 541 nsew
rlabel metal2 s 7818 14024 7926 14100 4 gnd
port 541 nsew
rlabel metal2 s 6570 16140 6678 16250 4 gnd
port 541 nsew
rlabel metal2 s 5802 1384 5910 1460 4 gnd
port 541 nsew
rlabel metal2 s 2826 15350 2934 15460 4 gnd
port 541 nsew
rlabel metal2 s 4554 21450 4662 21526 4 gnd
port 541 nsew
rlabel metal2 s 20778 1130 20886 1240 4 gnd
port 541 nsew
rlabel metal2 s 19050 23030 19158 23106 4 gnd
port 541 nsew
rlabel metal2 s 3306 24610 3414 24686 4 gnd
port 541 nsew
rlabel metal2 s 10794 11654 10902 11730 4 gnd
port 541 nsew
rlabel metal2 s 9546 4544 9654 4620 4 gnd
port 541 nsew
rlabel metal2 s 3306 1920 3414 2030 4 gnd
port 541 nsew
rlabel metal2 s 5802 10074 5910 10150 4 gnd
port 541 nsew
rlabel metal2 s 16554 20090 16662 20200 4 gnd
port 541 nsew
rlabel metal2 s 7050 12444 7158 12520 4 gnd
port 541 nsew
rlabel metal2 s 5802 3500 5910 3610 4 gnd
port 541 nsew
rlabel metal2 s 4074 910 4182 986 4 gnd
port 541 nsew
rlabel metal2 s 15786 9030 15894 9140 4 gnd
port 541 nsew
rlabel metal2 s 1578 7450 1686 7560 4 gnd
port 541 nsew
rlabel metal2 s 18282 13550 18390 13626 4 gnd
port 541 nsew
rlabel metal2 s 19530 12760 19638 12836 4 gnd
port 541 nsew
rlabel metal2 s 19530 5650 19638 5726 4 gnd
port 541 nsew
rlabel metal2 s 16554 13234 16662 13310 4 gnd
port 541 nsew
rlabel metal2 s 1578 5080 1686 5190 4 gnd
port 541 nsew
rlabel metal2 s 4074 13234 4182 13310 4 gnd
port 541 nsew
rlabel metal2 s 3306 12760 3414 12836 4 gnd
port 541 nsew
rlabel metal2 s 19050 22714 19158 22790 4 gnd
port 541 nsew
rlabel metal2 s 16554 7704 16662 7780 4 gnd
port 541 nsew
rlabel metal2 s 17802 340 17910 450 4 gnd
port 541 nsew
rlabel metal2 s 4554 19554 4662 19630 4 gnd
port 541 nsew
rlabel metal2 s 9546 120 9654 196 4 gnd
port 541 nsew
rlabel metal2 s 12042 2710 12150 2820 4 gnd
port 541 nsew
rlabel metal2 s 16554 4070 16662 4146 4 gnd
port 541 nsew
rlabel metal2 s 15306 23030 15414 23106 4 gnd
port 541 nsew
rlabel metal2 s 2826 10610 2934 10720 4 gnd
port 541 nsew
rlabel metal2 s 7050 15920 7158 15996 4 gnd
port 541 nsew
rlabel metal2 s 10314 18510 10422 18620 4 gnd
port 541 nsew
rlabel metal2 s 3306 17974 3414 18050 4 gnd
port 541 nsew
rlabel metal2 s 17802 21670 17910 21780 4 gnd
port 541 nsew
rlabel metal2 s 19050 20880 19158 20990 4 gnd
port 541 nsew
rlabel metal2 s 10794 340 10902 450 4 gnd
port 541 nsew
rlabel metal2 s 330 21670 438 21780 4 gnd
port 541 nsew
rlabel metal2 s 17034 5650 17142 5726 4 gnd
port 541 nsew
rlabel metal2 s 5322 11400 5430 11510 4 gnd
port 541 nsew
rlabel metal2 s 17802 20660 17910 20736 4 gnd
port 541 nsew
rlabel metal2 s 1578 10610 1686 10720 4 gnd
port 541 nsew
rlabel metal2 s 14538 15130 14646 15206 4 gnd
port 541 nsew
rlabel metal2 s 4074 12190 4182 12300 4 gnd
port 541 nsew
rlabel metal2 s 14538 11654 14646 11730 4 gnd
port 541 nsew
rlabel metal2 s 4074 19300 4182 19410 4 gnd
port 541 nsew
rlabel metal2 s 2058 6914 2166 6990 4 gnd
port 541 nsew
rlabel metal2 s 15306 14814 15414 14890 4 gnd
port 541 nsew
rlabel metal2 s 7818 13550 7926 13626 4 gnd
port 541 nsew
rlabel metal2 s 12810 10390 12918 10466 4 gnd
port 541 nsew
rlabel metal2 s 7050 14024 7158 14100 4 gnd
port 541 nsew
rlabel metal2 s 19050 8020 19158 8096 4 gnd
port 541 nsew
rlabel metal2 s 12810 16394 12918 16470 4 gnd
port 541 nsew
rlabel metal2 s 17034 25400 17142 25476 4 gnd
port 541 nsew
rlabel metal2 s 16554 2710 16662 2820 4 gnd
port 541 nsew
rlabel metal2 s 5322 16140 5430 16250 4 gnd
port 541 nsew
rlabel metal2 s 19050 4860 19158 4936 4 gnd
port 541 nsew
rlabel metal2 s 8298 6440 8406 6516 4 gnd
port 541 nsew
rlabel metal2 s 7818 16930 7926 17040 4 gnd
port 541 nsew
rlabel metal2 s 13290 11400 13398 11510 4 gnd
port 541 nsew
rlabel metal2 s 8298 17500 8406 17576 4 gnd
port 541 nsew
rlabel metal2 s 810 5334 918 5410 4 gnd
port 541 nsew
rlabel metal2 s 330 20090 438 20200 4 gnd
port 541 nsew
rlabel metal2 s 6570 6440 6678 6516 4 gnd
port 541 nsew
rlabel metal2 s 10314 1920 10422 2030 4 gnd
port 541 nsew
rlabel metal2 s 11562 340 11670 450 4 gnd
port 541 nsew
rlabel metal2 s 16554 9030 16662 9140 4 gnd
port 541 nsew
rlabel metal2 s 17034 594 17142 670 4 gnd
port 541 nsew
rlabel metal2 s 7050 3754 7158 3830 4 gnd
port 541 nsew
rlabel metal2 s 9546 18764 9654 18840 4 gnd
port 541 nsew
rlabel metal2 s 14538 24294 14646 24370 4 gnd
port 541 nsew
rlabel metal2 s 19050 14814 19158 14890 4 gnd
port 541 nsew
rlabel metal2 s 19530 21670 19638 21780 4 gnd
port 541 nsew
rlabel metal2 s 12810 17184 12918 17260 4 gnd
port 541 nsew
rlabel metal2 s 15306 6660 15414 6770 4 gnd
port 541 nsew
rlabel metal2 s 4074 10390 4182 10466 4 gnd
port 541 nsew
rlabel metal2 s 16554 23820 16662 23896 4 gnd
port 541 nsew
rlabel metal2 s 7050 14340 7158 14416 4 gnd
port 541 nsew
rlabel metal2 s 7050 13234 7158 13310 4 gnd
port 541 nsew
rlabel metal2 s 16554 1920 16662 2030 4 gnd
port 541 nsew
rlabel metal2 s 12042 8020 12150 8096 4 gnd
port 541 nsew
rlabel metal2 s 2058 340 2166 450 4 gnd
port 541 nsew
rlabel metal2 s 9546 19080 9654 19156 4 gnd
port 541 nsew
rlabel metal2 s 2826 17184 2934 17260 4 gnd
port 541 nsew
rlabel metal2 s 8298 23504 8406 23580 4 gnd
port 541 nsew
rlabel metal2 s 20298 19080 20406 19156 4 gnd
port 541 nsew
rlabel metal2 s 9546 13770 9654 13880 4 gnd
port 541 nsew
rlabel metal2 s 330 16394 438 16470 4 gnd
port 541 nsew
rlabel metal2 s 14058 5870 14166 5980 4 gnd
port 541 nsew
rlabel metal2 s 8298 19870 8406 19946 4 gnd
port 541 nsew
rlabel metal2 s 13290 14340 13398 14416 4 gnd
port 541 nsew
rlabel metal2 s 5802 15350 5910 15460 4 gnd
port 541 nsew
rlabel metal2 s 10314 6440 10422 6516 4 gnd
port 541 nsew
rlabel metal2 s 10794 15920 10902 15996 4 gnd
port 541 nsew
rlabel metal2 s 1578 4070 1686 4146 4 gnd
port 541 nsew
rlabel metal2 s 10314 24610 10422 24686 4 gnd
port 541 nsew
rlabel metal2 s 12042 13550 12150 13626 4 gnd
port 541 nsew
rlabel metal2 s 20778 20090 20886 20200 4 gnd
port 541 nsew
rlabel metal2 s 12810 13770 12918 13880 4 gnd
port 541 nsew
rlabel metal2 s 19050 17500 19158 17576 4 gnd
port 541 nsew
rlabel metal2 s 14538 21924 14646 22000 4 gnd
port 541 nsew
rlabel metal2 s 14058 12980 14166 13090 4 gnd
port 541 nsew
rlabel metal2 s 810 23504 918 23580 4 gnd
port 541 nsew
rlabel metal2 s 10314 12760 10422 12836 4 gnd
port 541 nsew
rlabel metal2 s 810 5080 918 5190 4 gnd
port 541 nsew
rlabel metal2 s 4074 16394 4182 16470 4 gnd
port 541 nsew
rlabel metal2 s 10314 24830 10422 24940 4 gnd
port 541 nsew
rlabel metal2 s 4554 19870 4662 19946 4 gnd
port 541 nsew
rlabel metal2 s 13290 14814 13398 14890 4 gnd
port 541 nsew
rlabel metal2 s 8298 16394 8406 16470 4 gnd
port 541 nsew
rlabel metal2 s 6570 21134 6678 21210 4 gnd
port 541 nsew
rlabel metal2 s 5802 19870 5910 19946 4 gnd
port 541 nsew
rlabel metal2 s 330 1384 438 1460 4 gnd
port 541 nsew
rlabel metal2 s 2826 10074 2934 10150 4 gnd
port 541 nsew
rlabel metal2 s 12042 340 12150 450 4 gnd
port 541 nsew
rlabel metal2 s 10314 22240 10422 22316 4 gnd
port 541 nsew
rlabel metal2 s 14058 5080 14166 5190 4 gnd
port 541 nsew
rlabel metal2 s 12810 17500 12918 17576 4 gnd
port 541 nsew
rlabel metal2 s 20298 7450 20406 7560 4 gnd
port 541 nsew
rlabel metal2 s 12810 20660 12918 20736 4 gnd
port 541 nsew
rlabel metal2 s 10314 7230 10422 7306 4 gnd
port 541 nsew
rlabel metal2 s 20298 8240 20406 8350 4 gnd
port 541 nsew
rlabel metal2 s 3306 8020 3414 8096 4 gnd
port 541 nsew
rlabel metal2 s 16554 19870 16662 19946 4 gnd
port 541 nsew
rlabel metal2 s 3306 24830 3414 24940 4 gnd
port 541 nsew
rlabel metal2 s 8298 20660 8406 20736 4 gnd
port 541 nsew
rlabel metal2 s 17802 18510 17910 18620 4 gnd
port 541 nsew
rlabel metal2 s 10314 11654 10422 11730 4 gnd
port 541 nsew
rlabel metal2 s 9546 16930 9654 17040 4 gnd
port 541 nsew
rlabel metal2 s 330 14340 438 14416 4 gnd
port 541 nsew
rlabel metal2 s 1578 13234 1686 13310 4 gnd
port 541 nsew
rlabel metal2 s 20298 13234 20406 13310 4 gnd
port 541 nsew
rlabel metal2 s 17034 18510 17142 18620 4 gnd
port 541 nsew
rlabel metal2 s 7818 19554 7926 19630 4 gnd
port 541 nsew
rlabel metal2 s 18282 6124 18390 6200 4 gnd
port 541 nsew
rlabel metal2 s 8298 22460 8406 22570 4 gnd
port 541 nsew
rlabel metal2 s 14058 7450 14166 7560 4 gnd
port 541 nsew
rlabel metal2 s 9066 15350 9174 15460 4 gnd
port 541 nsew
rlabel metal2 s 12810 1384 12918 1460 4 gnd
port 541 nsew
rlabel metal2 s 19050 594 19158 670 4 gnd
port 541 nsew
rlabel metal2 s 5802 25620 5910 25730 4 gnd
port 541 nsew
rlabel metal2 s 810 24830 918 24940 4 gnd
port 541 nsew
rlabel metal2 s 9066 4544 9174 4620 4 gnd
port 541 nsew
rlabel metal2 s 20778 15604 20886 15680 4 gnd
port 541 nsew
rlabel metal2 s 14538 20880 14646 20990 4 gnd
port 541 nsew
rlabel metal2 s 810 21134 918 21210 4 gnd
port 541 nsew
rlabel metal2 s 2058 18764 2166 18840 4 gnd
port 541 nsew
rlabel metal2 s 10794 5870 10902 5980 4 gnd
port 541 nsew
rlabel metal2 s 2058 594 2166 670 4 gnd
port 541 nsew
rlabel metal2 s 330 15604 438 15680 4 gnd
port 541 nsew
rlabel metal2 s 3306 16394 3414 16470 4 gnd
port 541 nsew
rlabel metal2 s 14538 340 14646 450 4 gnd
port 541 nsew
rlabel metal2 s 11562 22714 11670 22790 4 gnd
port 541 nsew
rlabel metal2 s 5322 21670 5430 21780 4 gnd
port 541 nsew
rlabel metal2 s 12042 910 12150 986 4 gnd
port 541 nsew
rlabel metal2 s 12042 23250 12150 23360 4 gnd
port 541 nsew
rlabel metal2 s 9546 3280 9654 3356 4 gnd
port 541 nsew
rlabel metal2 s 15786 9600 15894 9676 4 gnd
port 541 nsew
rlabel metal2 s 11562 2710 11670 2820 4 gnd
port 541 nsew
rlabel metal2 s 19530 594 19638 670 4 gnd
port 541 nsew
rlabel metal2 s 4554 7704 4662 7780 4 gnd
port 541 nsew
rlabel metal2 s 6570 24040 6678 24150 4 gnd
port 541 nsew
rlabel metal2 s 8298 16710 8406 16786 4 gnd
port 541 nsew
rlabel metal2 s 810 5650 918 5726 4 gnd
port 541 nsew
rlabel metal2 s 12042 15350 12150 15460 4 gnd
port 541 nsew
rlabel metal2 s 10314 19300 10422 19410 4 gnd
port 541 nsew
rlabel metal2 s 1578 19870 1686 19946 4 gnd
port 541 nsew
rlabel metal2 s 20778 25620 20886 25730 4 gnd
port 541 nsew
rlabel metal2 s 14538 4544 14646 4620 4 gnd
port 541 nsew
rlabel metal2 s 3306 23250 3414 23360 4 gnd
port 541 nsew
rlabel metal2 s 19050 11400 19158 11510 4 gnd
port 541 nsew
rlabel metal2 s 2058 13770 2166 13880 4 gnd
port 541 nsew
rlabel metal2 s 19050 25084 19158 25160 4 gnd
port 541 nsew
rlabel metal2 s 13290 25400 13398 25476 4 gnd
port 541 nsew
rlabel metal2 s 810 6440 918 6516 4 gnd
port 541 nsew
rlabel metal2 s 14058 594 14166 670 4 gnd
port 541 nsew
rlabel metal2 s 810 9030 918 9140 4 gnd
port 541 nsew
rlabel metal2 s 9066 20090 9174 20200 4 gnd
port 541 nsew
rlabel metal2 s 19050 14024 19158 14100 4 gnd
port 541 nsew
rlabel metal2 s 15306 5080 15414 5190 4 gnd
port 541 nsew
rlabel metal2 s 20298 16710 20406 16786 4 gnd
port 541 nsew
rlabel metal2 s 6570 12444 6678 12520 4 gnd
port 541 nsew
rlabel metal2 s 7050 6914 7158 6990 4 gnd
port 541 nsew
rlabel metal2 s 15786 21450 15894 21526 4 gnd
port 541 nsew
rlabel metal2 s 14538 7704 14646 7780 4 gnd
port 541 nsew
rlabel metal2 s 4074 4860 4182 4936 4 gnd
port 541 nsew
rlabel metal2 s 19050 20344 19158 20420 4 gnd
port 541 nsew
rlabel metal2 s 330 16930 438 17040 4 gnd
port 541 nsew
rlabel metal2 s 20778 21450 20886 21526 4 gnd
port 541 nsew
rlabel metal2 s 10794 17184 10902 17260 4 gnd
port 541 nsew
rlabel metal2 s 12042 23820 12150 23896 4 gnd
port 541 nsew
rlabel metal2 s 330 7450 438 7560 4 gnd
port 541 nsew
rlabel metal2 s 9546 8020 9654 8096 4 gnd
port 541 nsew
rlabel metal2 s 12810 9820 12918 9930 4 gnd
port 541 nsew
rlabel metal2 s 810 120 918 196 4 gnd
port 541 nsew
rlabel metal2 s 3306 2710 3414 2820 4 gnd
port 541 nsew
rlabel metal2 s 17034 11400 17142 11510 4 gnd
port 541 nsew
rlabel metal2 s 13290 17974 13398 18050 4 gnd
port 541 nsew
rlabel metal2 s 5802 1700 5910 1776 4 gnd
port 541 nsew
rlabel metal2 s 2826 4544 2934 4620 4 gnd
port 541 nsew
rlabel metal2 s 4074 15604 4182 15680 4 gnd
port 541 nsew
rlabel metal2 s 10794 22714 10902 22790 4 gnd
port 541 nsew
rlabel metal2 s 9066 20880 9174 20990 4 gnd
port 541 nsew
rlabel metal2 s 330 17184 438 17260 4 gnd
port 541 nsew
rlabel metal2 s 19530 340 19638 450 4 gnd
port 541 nsew
rlabel metal2 s 20778 10610 20886 10720 4 gnd
port 541 nsew
rlabel metal2 s 9066 9820 9174 9930 4 gnd
port 541 nsew
rlabel metal2 s 17802 22460 17910 22570 4 gnd
port 541 nsew
rlabel metal2 s 5802 24294 5910 24370 4 gnd
port 541 nsew
rlabel metal2 s 810 10390 918 10466 4 gnd
port 541 nsew
rlabel metal2 s 12810 8810 12918 8886 4 gnd
port 541 nsew
rlabel metal2 s 12042 10390 12150 10466 4 gnd
port 541 nsew
rlabel metal2 s 10314 2964 10422 3040 4 gnd
port 541 nsew
rlabel metal2 s 14058 13550 14166 13626 4 gnd
port 541 nsew
rlabel metal2 s 16554 25874 16662 25950 4 gnd
port 541 nsew
rlabel metal2 s 7818 11400 7926 11510 4 gnd
port 541 nsew
rlabel metal2 s 5322 11654 5430 11730 4 gnd
port 541 nsew
rlabel metal2 s 2826 23030 2934 23106 4 gnd
port 541 nsew
rlabel metal2 s 2826 13770 2934 13880 4 gnd
port 541 nsew
rlabel metal2 s 3306 4070 3414 4146 4 gnd
port 541 nsew
rlabel metal2 s 4554 23030 4662 23106 4 gnd
port 541 nsew
rlabel metal2 s 6570 16930 6678 17040 4 gnd
port 541 nsew
rlabel metal2 s 2058 8494 2166 8570 4 gnd
port 541 nsew
rlabel metal2 s 4074 21924 4182 22000 4 gnd
port 541 nsew
rlabel metal2 s 330 8810 438 8886 4 gnd
port 541 nsew
rlabel metal2 s 17802 18764 17910 18840 4 gnd
port 541 nsew
rlabel metal2 s 13290 25084 13398 25160 4 gnd
port 541 nsew
rlabel metal2 s 3306 10074 3414 10150 4 gnd
port 541 nsew
rlabel metal2 s 14058 20660 14166 20736 4 gnd
port 541 nsew
rlabel metal2 s 16554 24610 16662 24686 4 gnd
port 541 nsew
rlabel metal2 s 810 16710 918 16786 4 gnd
port 541 nsew
rlabel metal2 s 10314 20880 10422 20990 4 gnd
port 541 nsew
rlabel metal2 s 17802 2490 17910 2566 4 gnd
port 541 nsew
rlabel metal2 s 810 13234 918 13310 4 gnd
port 541 nsew
rlabel metal2 s 9066 8020 9174 8096 4 gnd
port 541 nsew
rlabel metal2 s 14058 10390 14166 10466 4 gnd
port 541 nsew
rlabel metal2 s 9066 21924 9174 22000 4 gnd
port 541 nsew
rlabel metal2 s 1578 16140 1686 16250 4 gnd
port 541 nsew
rlabel metal2 s 16554 20660 16662 20736 4 gnd
port 541 nsew
rlabel metal2 s 5322 25620 5430 25730 4 gnd
port 541 nsew
rlabel metal2 s 2826 910 2934 986 4 gnd
port 541 nsew
rlabel metal2 s 14058 15920 14166 15996 4 gnd
port 541 nsew
rlabel metal2 s 9546 25400 9654 25476 4 gnd
port 541 nsew
rlabel metal2 s 8298 4290 8406 4400 4 gnd
port 541 nsew
rlabel metal2 s 14538 14024 14646 14100 4 gnd
port 541 nsew
rlabel metal2 s 4074 25084 4182 25160 4 gnd
port 541 nsew
rlabel metal2 s 5802 22240 5910 22316 4 gnd
port 541 nsew
rlabel metal2 s 2058 13550 2166 13626 4 gnd
port 541 nsew
rlabel metal2 s 7818 14560 7926 14670 4 gnd
port 541 nsew
rlabel metal2 s 20778 2490 20886 2566 4 gnd
port 541 nsew
rlabel metal2 s 14058 6440 14166 6516 4 gnd
port 541 nsew
rlabel metal2 s 19530 9284 19638 9360 4 gnd
port 541 nsew
rlabel metal2 s 2058 6440 2166 6516 4 gnd
port 541 nsew
rlabel metal2 s 8298 3280 8406 3356 4 gnd
port 541 nsew
rlabel metal2 s 7050 14560 7158 14670 4 gnd
port 541 nsew
rlabel metal2 s 19050 15350 19158 15460 4 gnd
port 541 nsew
rlabel metal2 s 19050 17720 19158 17830 4 gnd
port 541 nsew
rlabel metal2 s 16554 910 16662 986 4 gnd
port 541 nsew
rlabel metal2 s 10314 11400 10422 11510 4 gnd
port 541 nsew
rlabel metal2 s 15306 8240 15414 8350 4 gnd
port 541 nsew
rlabel metal2 s 8298 16930 8406 17040 4 gnd
port 541 nsew
rlabel metal2 s 17034 13550 17142 13626 4 gnd
port 541 nsew
rlabel metal2 s 17034 340 17142 450 4 gnd
port 541 nsew
rlabel metal2 s 17034 10390 17142 10466 4 gnd
port 541 nsew
rlabel metal2 s 810 19300 918 19410 4 gnd
port 541 nsew
rlabel metal2 s 8298 9820 8406 9930 4 gnd
port 541 nsew
rlabel metal2 s 14538 23504 14646 23580 4 gnd
port 541 nsew
rlabel metal2 s 1578 18510 1686 18620 4 gnd
port 541 nsew
rlabel metal2 s 7050 20880 7158 20990 4 gnd
port 541 nsew
rlabel metal2 s 14058 6124 14166 6200 4 gnd
port 541 nsew
rlabel metal2 s 16554 21450 16662 21526 4 gnd
port 541 nsew
rlabel metal2 s 330 9284 438 9360 4 gnd
port 541 nsew
rlabel metal2 s 13290 3280 13398 3356 4 gnd
port 541 nsew
rlabel metal2 s 12810 24040 12918 24150 4 gnd
port 541 nsew
rlabel metal2 s 18282 23250 18390 23360 4 gnd
port 541 nsew
rlabel metal2 s 20778 18290 20886 18366 4 gnd
port 541 nsew
rlabel metal2 s 20298 21450 20406 21526 4 gnd
port 541 nsew
rlabel metal2 s 16554 9600 16662 9676 4 gnd
port 541 nsew
rlabel metal2 s 19050 17974 19158 18050 4 gnd
port 541 nsew
rlabel metal2 s 5802 1920 5910 2030 4 gnd
port 541 nsew
rlabel metal2 s 10794 11180 10902 11256 4 gnd
port 541 nsew
rlabel metal2 s 17034 3754 17142 3830 4 gnd
port 541 nsew
rlabel metal2 s 9066 1130 9174 1240 4 gnd
port 541 nsew
rlabel metal2 s 3306 6124 3414 6200 4 gnd
port 541 nsew
rlabel metal2 s 3306 10390 3414 10466 4 gnd
port 541 nsew
rlabel metal2 s 17034 4860 17142 4936 4 gnd
port 541 nsew
rlabel metal2 s 330 21450 438 21526 4 gnd
port 541 nsew
rlabel metal2 s 12810 3754 12918 3830 4 gnd
port 541 nsew
rlabel metal2 s 12042 4070 12150 4146 4 gnd
port 541 nsew
rlabel metal2 s 15306 11400 15414 11510 4 gnd
port 541 nsew
rlabel metal2 s 19530 16710 19638 16786 4 gnd
port 541 nsew
rlabel metal2 s 4554 4070 4662 4146 4 gnd
port 541 nsew
rlabel metal2 s 5802 5334 5910 5410 4 gnd
port 541 nsew
rlabel metal2 s 15786 22714 15894 22790 4 gnd
port 541 nsew
rlabel metal2 s 5322 8494 5430 8570 4 gnd
port 541 nsew
rlabel metal2 s 15786 20344 15894 20420 4 gnd
port 541 nsew
rlabel metal2 s 14058 18510 14166 18620 4 gnd
port 541 nsew
rlabel metal2 s 2058 12980 2166 13090 4 gnd
port 541 nsew
rlabel metal2 s 13290 340 13398 450 4 gnd
port 541 nsew
rlabel metal2 s 20778 18764 20886 18840 4 gnd
port 541 nsew
rlabel metal2 s 6570 12760 6678 12836 4 gnd
port 541 nsew
rlabel metal2 s 14538 2174 14646 2250 4 gnd
port 541 nsew
rlabel metal2 s 20298 25620 20406 25730 4 gnd
port 541 nsew
rlabel metal2 s 12042 22460 12150 22570 4 gnd
port 541 nsew
rlabel metal2 s 4074 24040 4182 24150 4 gnd
port 541 nsew
rlabel metal2 s 810 4544 918 4620 4 gnd
port 541 nsew
rlabel metal2 s 3306 5334 3414 5410 4 gnd
port 541 nsew
rlabel metal2 s 5322 6914 5430 6990 4 gnd
port 541 nsew
rlabel metal2 s 18282 20660 18390 20736 4 gnd
port 541 nsew
rlabel metal2 s 4074 9600 4182 9676 4 gnd
port 541 nsew
rlabel metal2 s 10314 10074 10422 10150 4 gnd
port 541 nsew
rlabel metal2 s 20298 12980 20406 13090 4 gnd
port 541 nsew
rlabel metal2 s 15786 4544 15894 4620 4 gnd
port 541 nsew
rlabel metal2 s 1578 6124 1686 6200 4 gnd
port 541 nsew
rlabel metal2 s 9546 16710 9654 16786 4 gnd
port 541 nsew
rlabel metal2 s 330 24830 438 24940 4 gnd
port 541 nsew
rlabel metal2 s 14058 14560 14166 14670 4 gnd
port 541 nsew
rlabel metal2 s 3306 15350 3414 15460 4 gnd
port 541 nsew
rlabel metal2 s 20298 10610 20406 10720 4 gnd
port 541 nsew
rlabel metal2 s 20298 12190 20406 12300 4 gnd
port 541 nsew
rlabel metal2 s 5802 12980 5910 13090 4 gnd
port 541 nsew
rlabel metal2 s 19530 8020 19638 8096 4 gnd
port 541 nsew
rlabel metal2 s 7818 18290 7926 18366 4 gnd
port 541 nsew
rlabel metal2 s 810 19080 918 19156 4 gnd
port 541 nsew
rlabel metal2 s 14058 25874 14166 25950 4 gnd
port 541 nsew
rlabel metal2 s 9066 20344 9174 20420 4 gnd
port 541 nsew
rlabel metal2 s 17802 4544 17910 4620 4 gnd
port 541 nsew
rlabel metal2 s 19530 19300 19638 19410 4 gnd
port 541 nsew
rlabel metal2 s 17034 6660 17142 6770 4 gnd
port 541 nsew
rlabel metal2 s 9066 19554 9174 19630 4 gnd
port 541 nsew
rlabel metal2 s 10794 10390 10902 10466 4 gnd
port 541 nsew
rlabel metal2 s 17802 594 17910 670 4 gnd
port 541 nsew
rlabel metal2 s 5802 20344 5910 20420 4 gnd
port 541 nsew
rlabel metal2 s 20298 17720 20406 17830 4 gnd
port 541 nsew
rlabel metal2 s 17802 10074 17910 10150 4 gnd
port 541 nsew
rlabel metal2 s 12042 11654 12150 11730 4 gnd
port 541 nsew
rlabel metal2 s 14058 21670 14166 21780 4 gnd
port 541 nsew
rlabel metal2 s 10794 19300 10902 19410 4 gnd
port 541 nsew
rlabel metal2 s 12042 18290 12150 18366 4 gnd
port 541 nsew
rlabel metal2 s 12810 7704 12918 7780 4 gnd
port 541 nsew
rlabel metal2 s 15786 7704 15894 7780 4 gnd
port 541 nsew
rlabel metal2 s 810 7230 918 7306 4 gnd
port 541 nsew
rlabel metal2 s 9066 17500 9174 17576 4 gnd
port 541 nsew
rlabel metal2 s 19530 14024 19638 14100 4 gnd
port 541 nsew
rlabel metal2 s 2826 10390 2934 10466 4 gnd
port 541 nsew
rlabel metal2 s 20298 2710 20406 2820 4 gnd
port 541 nsew
rlabel metal2 s 18282 25874 18390 25950 4 gnd
port 541 nsew
rlabel metal2 s 5802 25400 5910 25476 4 gnd
port 541 nsew
rlabel metal2 s 9546 2964 9654 3040 4 gnd
port 541 nsew
rlabel metal2 s 18282 2174 18390 2250 4 gnd
port 541 nsew
rlabel metal2 s 17034 2174 17142 2250 4 gnd
port 541 nsew
rlabel metal2 s 14538 17720 14646 17830 4 gnd
port 541 nsew
rlabel metal2 s 10794 7230 10902 7306 4 gnd
port 541 nsew
rlabel metal2 s 8298 20090 8406 20200 4 gnd
port 541 nsew
rlabel metal2 s 2058 23504 2166 23580 4 gnd
port 541 nsew
rlabel metal2 s 10314 8810 10422 8886 4 gnd
port 541 nsew
rlabel metal2 s 16554 15920 16662 15996 4 gnd
port 541 nsew
rlabel metal2 s 14538 5080 14646 5190 4 gnd
port 541 nsew
rlabel metal2 s 16554 18510 16662 18620 4 gnd
port 541 nsew
rlabel metal2 s 12042 14814 12150 14890 4 gnd
port 541 nsew
rlabel metal2 s 14538 22240 14646 22316 4 gnd
port 541 nsew
rlabel metal2 s 16554 22240 16662 22316 4 gnd
port 541 nsew
rlabel metal2 s 2826 7230 2934 7306 4 gnd
port 541 nsew
rlabel metal2 s 7818 6660 7926 6770 4 gnd
port 541 nsew
rlabel metal2 s 20298 11400 20406 11510 4 gnd
port 541 nsew
rlabel metal2 s 15306 1384 15414 1460 4 gnd
port 541 nsew
rlabel metal2 s 14538 3754 14646 3830 4 gnd
port 541 nsew
rlabel metal2 s 14058 6914 14166 6990 4 gnd
port 541 nsew
rlabel metal2 s 5322 15130 5430 15206 4 gnd
port 541 nsew
rlabel metal2 s 8298 19554 8406 19630 4 gnd
port 541 nsew
rlabel metal2 s 20778 594 20886 670 4 gnd
port 541 nsew
rlabel metal2 s 5322 17500 5430 17576 4 gnd
port 541 nsew
rlabel metal2 s 810 18290 918 18366 4 gnd
port 541 nsew
rlabel metal2 s 810 21924 918 22000 4 gnd
port 541 nsew
rlabel metal2 s 17802 11970 17910 12046 4 gnd
port 541 nsew
rlabel metal2 s 17034 12190 17142 12300 4 gnd
port 541 nsew
rlabel metal2 s 9066 22240 9174 22316 4 gnd
port 541 nsew
rlabel metal2 s 9066 16394 9174 16470 4 gnd
port 541 nsew
rlabel metal2 s 14058 25620 14166 25730 4 gnd
port 541 nsew
rlabel metal2 s 14058 6660 14166 6770 4 gnd
port 541 nsew
rlabel metal2 s 10314 23250 10422 23360 4 gnd
port 541 nsew
rlabel metal2 s 17802 4290 17910 4400 4 gnd
port 541 nsew
rlabel metal2 s 9546 17184 9654 17260 4 gnd
port 541 nsew
rlabel metal2 s 2826 6660 2934 6770 4 gnd
port 541 nsew
rlabel metal2 s 16554 10610 16662 10720 4 gnd
port 541 nsew
rlabel metal2 s 11562 594 11670 670 4 gnd
port 541 nsew
rlabel metal2 s 11562 5870 11670 5980 4 gnd
port 541 nsew
rlabel metal2 s 5802 9030 5910 9140 4 gnd
port 541 nsew
rlabel metal2 s 2826 7450 2934 7560 4 gnd
port 541 nsew
rlabel metal2 s 20298 13550 20406 13626 4 gnd
port 541 nsew
rlabel metal2 s 9066 15920 9174 15996 4 gnd
port 541 nsew
rlabel metal2 s 7050 20660 7158 20736 4 gnd
port 541 nsew
rlabel metal2 s 9066 19300 9174 19410 4 gnd
port 541 nsew
rlabel metal2 s 810 15130 918 15206 4 gnd
port 541 nsew
rlabel metal2 s 5802 16930 5910 17040 4 gnd
port 541 nsew
rlabel metal2 s 3306 7230 3414 7306 4 gnd
port 541 nsew
rlabel metal2 s 4074 24830 4182 24940 4 gnd
port 541 nsew
rlabel metal2 s 6570 18290 6678 18366 4 gnd
port 541 nsew
rlabel metal2 s 15786 14560 15894 14670 4 gnd
port 541 nsew
rlabel metal2 s 13290 2174 13398 2250 4 gnd
port 541 nsew
rlabel metal2 s 2826 4860 2934 4936 4 gnd
port 541 nsew
rlabel metal2 s 15786 19554 15894 19630 4 gnd
port 541 nsew
rlabel metal2 s 2058 22714 2166 22790 4 gnd
port 541 nsew
rlabel metal2 s 4554 2964 4662 3040 4 gnd
port 541 nsew
rlabel metal2 s 7050 8020 7158 8096 4 gnd
port 541 nsew
rlabel metal2 s 14058 4290 14166 4400 4 gnd
port 541 nsew
rlabel metal2 s 9066 16710 9174 16786 4 gnd
port 541 nsew
rlabel metal2 s 15786 23820 15894 23896 4 gnd
port 541 nsew
rlabel metal2 s 12042 13770 12150 13880 4 gnd
port 541 nsew
rlabel metal2 s 8298 120 8406 196 4 gnd
port 541 nsew
rlabel metal2 s 19050 23820 19158 23896 4 gnd
port 541 nsew
rlabel metal2 s 6570 6660 6678 6770 4 gnd
port 541 nsew
rlabel metal2 s 12810 22460 12918 22570 4 gnd
port 541 nsew
rlabel metal2 s 16554 5650 16662 5726 4 gnd
port 541 nsew
rlabel metal2 s 14538 6440 14646 6516 4 gnd
port 541 nsew
rlabel metal2 s 14538 24040 14646 24150 4 gnd
port 541 nsew
rlabel metal2 s 20298 15920 20406 15996 4 gnd
port 541 nsew
rlabel metal2 s 9546 15920 9654 15996 4 gnd
port 541 nsew
rlabel metal2 s 12042 8810 12150 8886 4 gnd
port 541 nsew
rlabel metal2 s 17034 11180 17142 11256 4 gnd
port 541 nsew
rlabel metal2 s 7818 15350 7926 15460 4 gnd
port 541 nsew
rlabel metal2 s 7818 9820 7926 9930 4 gnd
port 541 nsew
rlabel metal2 s 14058 24830 14166 24940 4 gnd
port 541 nsew
rlabel metal2 s 8298 6914 8406 6990 4 gnd
port 541 nsew
rlabel metal2 s 4554 12980 4662 13090 4 gnd
port 541 nsew
rlabel metal2 s 15786 2710 15894 2820 4 gnd
port 541 nsew
rlabel metal2 s 4554 21924 4662 22000 4 gnd
port 541 nsew
rlabel metal2 s 6570 20090 6678 20200 4 gnd
port 541 nsew
rlabel metal2 s 16554 12980 16662 13090 4 gnd
port 541 nsew
rlabel metal2 s 8298 1920 8406 2030 4 gnd
port 541 nsew
rlabel metal2 s 5802 16710 5910 16786 4 gnd
port 541 nsew
rlabel metal2 s 17034 23030 17142 23106 4 gnd
port 541 nsew
rlabel metal2 s 12042 11180 12150 11256 4 gnd
port 541 nsew
rlabel metal2 s 5322 6660 5430 6770 4 gnd
port 541 nsew
rlabel metal2 s 8298 340 8406 450 4 gnd
port 541 nsew
rlabel metal2 s 9066 7704 9174 7780 4 gnd
port 541 nsew
rlabel metal2 s 3306 23504 3414 23580 4 gnd
port 541 nsew
rlabel metal2 s 14058 22460 14166 22570 4 gnd
port 541 nsew
rlabel metal2 s 9066 4070 9174 4146 4 gnd
port 541 nsew
rlabel metal2 s 14538 17500 14646 17576 4 gnd
port 541 nsew
rlabel metal2 s 15306 20344 15414 20420 4 gnd
port 541 nsew
rlabel metal2 s 4554 23250 4662 23360 4 gnd
port 541 nsew
rlabel metal2 s 2058 4070 2166 4146 4 gnd
port 541 nsew
rlabel metal2 s 16554 9284 16662 9360 4 gnd
port 541 nsew
rlabel metal2 s 9546 594 9654 670 4 gnd
port 541 nsew
rlabel metal2 s 20298 4544 20406 4620 4 gnd
port 541 nsew
rlabel metal2 s 17802 22714 17910 22790 4 gnd
port 541 nsew
rlabel metal2 s 2058 23820 2166 23896 4 gnd
port 541 nsew
rlabel metal2 s 7818 1920 7926 2030 4 gnd
port 541 nsew
rlabel metal2 s 10314 13550 10422 13626 4 gnd
port 541 nsew
rlabel metal2 s 2826 18764 2934 18840 4 gnd
port 541 nsew
rlabel metal2 s 4074 14024 4182 14100 4 gnd
port 541 nsew
rlabel metal2 s 13290 21450 13398 21526 4 gnd
port 541 nsew
rlabel metal2 s 18282 1384 18390 1460 4 gnd
port 541 nsew
rlabel metal2 s 14058 15130 14166 15206 4 gnd
port 541 nsew
rlabel metal2 s 20778 1920 20886 2030 4 gnd
port 541 nsew
rlabel metal2 s 15786 2490 15894 2566 4 gnd
port 541 nsew
rlabel metal2 s 810 340 918 450 4 gnd
port 541 nsew
rlabel metal2 s 15306 12760 15414 12836 4 gnd
port 541 nsew
rlabel metal2 s 13290 910 13398 986 4 gnd
port 541 nsew
rlabel metal2 s 4554 1920 4662 2030 4 gnd
port 541 nsew
rlabel metal2 s 9546 20344 9654 20420 4 gnd
port 541 nsew
rlabel metal2 s 10314 16930 10422 17040 4 gnd
port 541 nsew
rlabel metal2 s 15306 12980 15414 13090 4 gnd
port 541 nsew
rlabel metal2 s 12810 8020 12918 8096 4 gnd
port 541 nsew
rlabel metal2 s 7050 2964 7158 3040 4 gnd
port 541 nsew
rlabel metal2 s 1578 24294 1686 24370 4 gnd
port 541 nsew
rlabel metal2 s 11562 2174 11670 2250 4 gnd
port 541 nsew
rlabel metal2 s 3306 12980 3414 13090 4 gnd
port 541 nsew
rlabel metal2 s 5802 18764 5910 18840 4 gnd
port 541 nsew
rlabel metal2 s 1578 10390 1686 10466 4 gnd
port 541 nsew
rlabel metal2 s 20298 120 20406 196 4 gnd
port 541 nsew
rlabel metal2 s 13290 17184 13398 17260 4 gnd
port 541 nsew
rlabel metal2 s 5802 9820 5910 9930 4 gnd
port 541 nsew
rlabel metal2 s 6570 7450 6678 7560 4 gnd
port 541 nsew
rlabel metal2 s 7050 8240 7158 8350 4 gnd
port 541 nsew
rlabel metal2 s 11562 1700 11670 1776 4 gnd
port 541 nsew
rlabel metal2 s 17802 1384 17910 1460 4 gnd
port 541 nsew
rlabel metal2 s 10794 24610 10902 24686 4 gnd
port 541 nsew
rlabel metal2 s 4554 4544 4662 4620 4 gnd
port 541 nsew
rlabel metal2 s 5322 2490 5430 2566 4 gnd
port 541 nsew
rlabel metal2 s 9066 12760 9174 12836 4 gnd
port 541 nsew
rlabel metal2 s 5322 11970 5430 12046 4 gnd
port 541 nsew
rlabel metal2 s 7050 25400 7158 25476 4 gnd
port 541 nsew
rlabel metal2 s 14058 13234 14166 13310 4 gnd
port 541 nsew
rlabel metal2 s 7050 24830 7158 24940 4 gnd
port 541 nsew
rlabel metal2 s 14058 8810 14166 8886 4 gnd
port 541 nsew
rlabel metal2 s 8298 22240 8406 22316 4 gnd
port 541 nsew
rlabel metal2 s 6570 25620 6678 25730 4 gnd
port 541 nsew
rlabel metal2 s 10314 5650 10422 5726 4 gnd
port 541 nsew
rlabel metal2 s 3306 19554 3414 19630 4 gnd
port 541 nsew
rlabel metal2 s 2058 910 2166 986 4 gnd
port 541 nsew
rlabel metal2 s 17034 17974 17142 18050 4 gnd
port 541 nsew
rlabel metal2 s 7050 9820 7158 9930 4 gnd
port 541 nsew
rlabel metal2 s 6570 4544 6678 4620 4 gnd
port 541 nsew
rlabel metal2 s 19050 4544 19158 4620 4 gnd
port 541 nsew
rlabel metal2 s 2826 15604 2934 15680 4 gnd
port 541 nsew
rlabel metal2 s 14538 10610 14646 10720 4 gnd
port 541 nsew
rlabel metal2 s 7818 6440 7926 6516 4 gnd
port 541 nsew
rlabel metal2 s 3306 1130 3414 1240 4 gnd
port 541 nsew
rlabel metal2 s 12042 7704 12150 7780 4 gnd
port 541 nsew
rlabel metal2 s 14538 3500 14646 3610 4 gnd
port 541 nsew
rlabel metal2 s 19050 3754 19158 3830 4 gnd
port 541 nsew
rlabel metal2 s 19530 5870 19638 5980 4 gnd
port 541 nsew
rlabel metal2 s 8298 910 8406 986 4 gnd
port 541 nsew
rlabel metal2 s 13290 12760 13398 12836 4 gnd
port 541 nsew
rlabel metal2 s 17802 10390 17910 10466 4 gnd
port 541 nsew
rlabel metal2 s 15306 2964 15414 3040 4 gnd
port 541 nsew
rlabel metal2 s 19050 25400 19158 25476 4 gnd
port 541 nsew
rlabel metal2 s 5802 13770 5910 13880 4 gnd
port 541 nsew
rlabel metal2 s 12810 6660 12918 6770 4 gnd
port 541 nsew
rlabel metal2 s 15786 19080 15894 19156 4 gnd
port 541 nsew
rlabel metal2 s 5802 2174 5910 2250 4 gnd
port 541 nsew
rlabel metal2 s 4554 10074 4662 10150 4 gnd
port 541 nsew
rlabel metal2 s 11562 6660 11670 6770 4 gnd
port 541 nsew
rlabel metal2 s 19530 24294 19638 24370 4 gnd
port 541 nsew
rlabel metal2 s 18282 10610 18390 10720 4 gnd
port 541 nsew
rlabel metal2 s 2058 15350 2166 15460 4 gnd
port 541 nsew
rlabel metal2 s 20778 10390 20886 10466 4 gnd
port 541 nsew
rlabel metal2 s 15786 340 15894 450 4 gnd
port 541 nsew
rlabel metal2 s 7818 2964 7926 3040 4 gnd
port 541 nsew
rlabel metal2 s 8298 24294 8406 24370 4 gnd
port 541 nsew
rlabel metal2 s 10314 6124 10422 6200 4 gnd
port 541 nsew
rlabel metal2 s 1578 1384 1686 1460 4 gnd
port 541 nsew
rlabel metal2 s 9066 9284 9174 9360 4 gnd
port 541 nsew
rlabel metal2 s 1578 25084 1686 25160 4 gnd
port 541 nsew
rlabel metal2 s 4554 6124 4662 6200 4 gnd
port 541 nsew
rlabel metal2 s 2058 10074 2166 10150 4 gnd
port 541 nsew
rlabel metal2 s 17802 6914 17910 6990 4 gnd
port 541 nsew
rlabel metal2 s 16554 9820 16662 9930 4 gnd
port 541 nsew
rlabel metal2 s 19530 18290 19638 18366 4 gnd
port 541 nsew
rlabel metal2 s 2058 19080 2166 19156 4 gnd
port 541 nsew
rlabel metal2 s 5802 9600 5910 9676 4 gnd
port 541 nsew
rlabel metal2 s 330 24610 438 24686 4 gnd
port 541 nsew
rlabel metal2 s 18282 16394 18390 16470 4 gnd
port 541 nsew
rlabel metal2 s 19050 10864 19158 10940 4 gnd
port 541 nsew
rlabel metal2 s 2826 15130 2934 15206 4 gnd
port 541 nsew
rlabel metal2 s 9546 21450 9654 21526 4 gnd
port 541 nsew
rlabel metal2 s 810 4290 918 4400 4 gnd
port 541 nsew
rlabel metal2 s 1578 23030 1686 23106 4 gnd
port 541 nsew
rlabel metal2 s 1578 4860 1686 4936 4 gnd
port 541 nsew
rlabel metal2 s 17802 14024 17910 14100 4 gnd
port 541 nsew
rlabel metal2 s 5802 17974 5910 18050 4 gnd
port 541 nsew
rlabel metal2 s 10314 19870 10422 19946 4 gnd
port 541 nsew
rlabel metal2 s 4074 120 4182 196 4 gnd
port 541 nsew
rlabel metal2 s 19050 12444 19158 12520 4 gnd
port 541 nsew
rlabel metal2 s 16554 1384 16662 1460 4 gnd
port 541 nsew
rlabel metal2 s 17034 3500 17142 3610 4 gnd
port 541 nsew
rlabel metal2 s 12042 19554 12150 19630 4 gnd
port 541 nsew
rlabel metal2 s 13290 9030 13398 9140 4 gnd
port 541 nsew
rlabel metal2 s 19530 22714 19638 22790 4 gnd
port 541 nsew
rlabel metal2 s 14538 24610 14646 24686 4 gnd
port 541 nsew
rlabel metal2 s 3306 10610 3414 10720 4 gnd
port 541 nsew
rlabel metal2 s 4554 25084 4662 25160 4 gnd
port 541 nsew
rlabel metal2 s 7050 16140 7158 16250 4 gnd
port 541 nsew
rlabel metal2 s 17802 20880 17910 20990 4 gnd
port 541 nsew
rlabel metal2 s 5322 20090 5430 20200 4 gnd
port 541 nsew
rlabel metal2 s 14058 16710 14166 16786 4 gnd
port 541 nsew
rlabel metal2 s 6570 5334 6678 5410 4 gnd
port 541 nsew
rlabel metal2 s 18282 1920 18390 2030 4 gnd
port 541 nsew
rlabel metal2 s 15306 120 15414 196 4 gnd
port 541 nsew
rlabel metal2 s 2058 14560 2166 14670 4 gnd
port 541 nsew
rlabel metal2 s 17802 25620 17910 25730 4 gnd
port 541 nsew
rlabel metal2 s 2826 17720 2934 17830 4 gnd
port 541 nsew
rlabel metal2 s 16554 24830 16662 24940 4 gnd
port 541 nsew
rlabel metal2 s 4554 6914 4662 6990 4 gnd
port 541 nsew
rlabel metal2 s 19530 19080 19638 19156 4 gnd
port 541 nsew
rlabel metal2 s 10794 5650 10902 5726 4 gnd
port 541 nsew
rlabel metal2 s 14538 3280 14646 3356 4 gnd
port 541 nsew
rlabel metal2 s 15306 19300 15414 19410 4 gnd
port 541 nsew
rlabel metal2 s 14538 7230 14646 7306 4 gnd
port 541 nsew
rlabel metal2 s 19050 10610 19158 10720 4 gnd
port 541 nsew
rlabel metal2 s 810 3500 918 3610 4 gnd
port 541 nsew
rlabel metal2 s 19530 20880 19638 20990 4 gnd
port 541 nsew
rlabel metal2 s 8298 23250 8406 23360 4 gnd
port 541 nsew
rlabel metal2 s 1578 22460 1686 22570 4 gnd
port 541 nsew
rlabel metal2 s 3306 14560 3414 14670 4 gnd
port 541 nsew
rlabel metal2 s 12042 5870 12150 5980 4 gnd
port 541 nsew
rlabel metal2 s 4554 23504 4662 23580 4 gnd
port 541 nsew
rlabel metal2 s 17034 25084 17142 25160 4 gnd
port 541 nsew
rlabel metal2 s 12810 10074 12918 10150 4 gnd
port 541 nsew
rlabel metal2 s 6570 1700 6678 1776 4 gnd
port 541 nsew
rlabel metal2 s 13290 25620 13398 25730 4 gnd
port 541 nsew
rlabel metal2 s 12810 23250 12918 23360 4 gnd
port 541 nsew
rlabel metal2 s 2058 8020 2166 8096 4 gnd
port 541 nsew
rlabel metal2 s 14058 23820 14166 23896 4 gnd
port 541 nsew
rlabel metal2 s 7050 12190 7158 12300 4 gnd
port 541 nsew
rlabel metal2 s 8298 15350 8406 15460 4 gnd
port 541 nsew
rlabel metal2 s 10314 14560 10422 14670 4 gnd
port 541 nsew
rlabel metal2 s 2826 20344 2934 20420 4 gnd
port 541 nsew
rlabel metal2 s 810 20880 918 20990 4 gnd
port 541 nsew
rlabel metal2 s 15786 16394 15894 16470 4 gnd
port 541 nsew
rlabel metal2 s 11562 11654 11670 11730 4 gnd
port 541 nsew
rlabel metal2 s 3306 5080 3414 5190 4 gnd
port 541 nsew
rlabel metal2 s 4554 5334 4662 5410 4 gnd
port 541 nsew
rlabel metal2 s 17034 2964 17142 3040 4 gnd
port 541 nsew
rlabel metal2 s 12042 8494 12150 8570 4 gnd
port 541 nsew
rlabel metal2 s 2826 5650 2934 5726 4 gnd
port 541 nsew
rlabel metal2 s 19050 20660 19158 20736 4 gnd
port 541 nsew
rlabel metal2 s 4074 23820 4182 23896 4 gnd
port 541 nsew
rlabel metal2 s 19050 19080 19158 19156 4 gnd
port 541 nsew
rlabel metal2 s 7050 18510 7158 18620 4 gnd
port 541 nsew
rlabel metal2 s 20778 11180 20886 11256 4 gnd
port 541 nsew
rlabel metal2 s 7050 15130 7158 15206 4 gnd
port 541 nsew
rlabel metal2 s 19530 16930 19638 17040 4 gnd
port 541 nsew
rlabel metal2 s 20778 10864 20886 10940 4 gnd
port 541 nsew
rlabel metal2 s 1578 22240 1686 22316 4 gnd
port 541 nsew
rlabel metal2 s 5802 17720 5910 17830 4 gnd
port 541 nsew
rlabel metal2 s 10314 12980 10422 13090 4 gnd
port 541 nsew
rlabel metal2 s 2826 3500 2934 3610 4 gnd
port 541 nsew
rlabel metal2 s 10314 25400 10422 25476 4 gnd
port 541 nsew
rlabel metal2 s 9066 14814 9174 14890 4 gnd
port 541 nsew
rlabel metal2 s 10794 25084 10902 25160 4 gnd
port 541 nsew
rlabel metal2 s 4074 22240 4182 22316 4 gnd
port 541 nsew
rlabel metal2 s 16554 8810 16662 8886 4 gnd
port 541 nsew
rlabel metal2 s 5322 20344 5430 20420 4 gnd
port 541 nsew
rlabel metal2 s 7818 11654 7926 11730 4 gnd
port 541 nsew
rlabel metal2 s 12810 12190 12918 12300 4 gnd
port 541 nsew
rlabel metal2 s 12810 5334 12918 5410 4 gnd
port 541 nsew
rlabel metal2 s 14058 19080 14166 19156 4 gnd
port 541 nsew
rlabel metal2 s 3306 14340 3414 14416 4 gnd
port 541 nsew
rlabel metal2 s 20778 8240 20886 8350 4 gnd
port 541 nsew
rlabel metal2 s 14058 16140 14166 16250 4 gnd
port 541 nsew
rlabel metal2 s 9066 2174 9174 2250 4 gnd
port 541 nsew
rlabel metal2 s 5802 17500 5910 17576 4 gnd
port 541 nsew
rlabel metal2 s 14538 10864 14646 10940 4 gnd
port 541 nsew
rlabel metal2 s 7818 5334 7926 5410 4 gnd
port 541 nsew
rlabel metal2 s 13290 7230 13398 7306 4 gnd
port 541 nsew
rlabel metal2 s 2826 1920 2934 2030 4 gnd
port 541 nsew
rlabel metal2 s 17802 910 17910 986 4 gnd
port 541 nsew
rlabel metal2 s 16554 17720 16662 17830 4 gnd
port 541 nsew
rlabel metal2 s 3306 25400 3414 25476 4 gnd
port 541 nsew
rlabel metal2 s 15306 16930 15414 17040 4 gnd
port 541 nsew
rlabel metal2 s 13290 10864 13398 10940 4 gnd
port 541 nsew
rlabel metal2 s 2826 18290 2934 18366 4 gnd
port 541 nsew
rlabel metal2 s 14058 1700 14166 1776 4 gnd
port 541 nsew
rlabel metal2 s 2826 1700 2934 1776 4 gnd
port 541 nsew
rlabel metal2 s 19050 910 19158 986 4 gnd
port 541 nsew
rlabel metal2 s 7818 20344 7926 20420 4 gnd
port 541 nsew
rlabel metal2 s 12810 4070 12918 4146 4 gnd
port 541 nsew
rlabel metal2 s 330 5080 438 5190 4 gnd
port 541 nsew
rlabel metal2 s 10314 5080 10422 5190 4 gnd
port 541 nsew
rlabel metal2 s 16554 8020 16662 8096 4 gnd
port 541 nsew
rlabel metal2 s 330 21134 438 21210 4 gnd
port 541 nsew
rlabel metal2 s 20298 19870 20406 19946 4 gnd
port 541 nsew
rlabel metal2 s 12042 13234 12150 13310 4 gnd
port 541 nsew
rlabel metal2 s 7050 16710 7158 16786 4 gnd
port 541 nsew
rlabel metal2 s 4074 3280 4182 3356 4 gnd
port 541 nsew
rlabel metal2 s 5322 7704 5430 7780 4 gnd
port 541 nsew
rlabel metal2 s 13290 11970 13398 12046 4 gnd
port 541 nsew
rlabel metal2 s 9066 4290 9174 4400 4 gnd
port 541 nsew
rlabel metal2 s 9546 14340 9654 14416 4 gnd
port 541 nsew
rlabel metal2 s 18282 23504 18390 23580 4 gnd
port 541 nsew
rlabel metal2 s 10794 9820 10902 9930 4 gnd
port 541 nsew
rlabel metal2 s 19530 9600 19638 9676 4 gnd
port 541 nsew
rlabel metal2 s 18282 5870 18390 5980 4 gnd
port 541 nsew
rlabel metal2 s 15306 21134 15414 21210 4 gnd
port 541 nsew
rlabel metal2 s 18282 12190 18390 12300 4 gnd
port 541 nsew
rlabel metal2 s 16554 15350 16662 15460 4 gnd
port 541 nsew
rlabel metal2 s 14538 25874 14646 25950 4 gnd
port 541 nsew
rlabel metal2 s 9546 25874 9654 25950 4 gnd
port 541 nsew
rlabel metal2 s 15786 11400 15894 11510 4 gnd
port 541 nsew
rlabel metal2 s 5322 594 5430 670 4 gnd
port 541 nsew
rlabel metal2 s 14058 24040 14166 24150 4 gnd
port 541 nsew
rlabel metal2 s 13290 14560 13398 14670 4 gnd
port 541 nsew
rlabel metal2 s 5322 18290 5430 18366 4 gnd
port 541 nsew
rlabel metal2 s 12042 2174 12150 2250 4 gnd
port 541 nsew
rlabel metal2 s 11562 20344 11670 20420 4 gnd
port 541 nsew
rlabel metal2 s 4074 17500 4182 17576 4 gnd
port 541 nsew
rlabel metal2 s 18282 2490 18390 2566 4 gnd
port 541 nsew
rlabel metal2 s 6570 15350 6678 15460 4 gnd
port 541 nsew
rlabel metal2 s 9546 9820 9654 9930 4 gnd
port 541 nsew
rlabel metal2 s 8298 24040 8406 24150 4 gnd
port 541 nsew
rlabel metal2 s 14058 17720 14166 17830 4 gnd
port 541 nsew
rlabel metal2 s 6570 23250 6678 23360 4 gnd
port 541 nsew
rlabel metal2 s 1578 120 1686 196 4 gnd
port 541 nsew
rlabel metal2 s 18282 21670 18390 21780 4 gnd
port 541 nsew
rlabel metal2 s 19050 17184 19158 17260 4 gnd
port 541 nsew
rlabel metal2 s 19050 6660 19158 6770 4 gnd
port 541 nsew
rlabel metal2 s 5322 1920 5430 2030 4 gnd
port 541 nsew
rlabel metal2 s 10314 7704 10422 7780 4 gnd
port 541 nsew
rlabel metal2 s 2058 22460 2166 22570 4 gnd
port 541 nsew
rlabel metal2 s 17034 11654 17142 11730 4 gnd
port 541 nsew
rlabel metal2 s 4074 15350 4182 15460 4 gnd
port 541 nsew
rlabel metal2 s 2826 22240 2934 22316 4 gnd
port 541 nsew
rlabel metal2 s 15306 23250 15414 23360 4 gnd
port 541 nsew
rlabel metal2 s 4074 5080 4182 5190 4 gnd
port 541 nsew
rlabel metal2 s 12042 12760 12150 12836 4 gnd
port 541 nsew
rlabel metal2 s 17034 1130 17142 1240 4 gnd
port 541 nsew
rlabel metal2 s 17802 12980 17910 13090 4 gnd
port 541 nsew
rlabel metal2 s 8298 2490 8406 2566 4 gnd
port 541 nsew
rlabel metal2 s 14058 18764 14166 18840 4 gnd
port 541 nsew
rlabel metal2 s 20778 23504 20886 23580 4 gnd
port 541 nsew
rlabel metal2 s 8298 10610 8406 10720 4 gnd
port 541 nsew
rlabel metal2 s 7818 12760 7926 12836 4 gnd
port 541 nsew
rlabel metal2 s 15306 11970 15414 12046 4 gnd
port 541 nsew
rlabel metal2 s 10314 25874 10422 25950 4 gnd
port 541 nsew
rlabel metal2 s 17802 16710 17910 16786 4 gnd
port 541 nsew
rlabel metal2 s 1578 9600 1686 9676 4 gnd
port 541 nsew
rlabel metal2 s 18282 19300 18390 19410 4 gnd
port 541 nsew
rlabel metal2 s 12042 25620 12150 25730 4 gnd
port 541 nsew
rlabel metal2 s 330 19300 438 19410 4 gnd
port 541 nsew
rlabel metal2 s 17802 11654 17910 11730 4 gnd
port 541 nsew
rlabel metal2 s 15306 594 15414 670 4 gnd
port 541 nsew
rlabel metal2 s 13290 18764 13398 18840 4 gnd
port 541 nsew
rlabel metal2 s 19050 4070 19158 4146 4 gnd
port 541 nsew
rlabel metal2 s 8298 7450 8406 7560 4 gnd
port 541 nsew
rlabel metal2 s 16554 6124 16662 6200 4 gnd
port 541 nsew
rlabel metal2 s 9546 23030 9654 23106 4 gnd
port 541 nsew
rlabel metal2 s 13290 10074 13398 10150 4 gnd
port 541 nsew
rlabel metal2 s 14058 25400 14166 25476 4 gnd
port 541 nsew
rlabel metal2 s 12810 24610 12918 24686 4 gnd
port 541 nsew
rlabel metal2 s 2058 7450 2166 7560 4 gnd
port 541 nsew
rlabel metal2 s 6570 16710 6678 16786 4 gnd
port 541 nsew
rlabel metal2 s 7818 17500 7926 17576 4 gnd
port 541 nsew
rlabel metal2 s 14058 16394 14166 16470 4 gnd
port 541 nsew
rlabel metal2 s 14058 24294 14166 24370 4 gnd
port 541 nsew
rlabel metal2 s 19050 5080 19158 5190 4 gnd
port 541 nsew
rlabel metal2 s 3306 9284 3414 9360 4 gnd
port 541 nsew
rlabel metal2 s 17802 20090 17910 20200 4 gnd
port 541 nsew
rlabel metal2 s 3306 2964 3414 3040 4 gnd
port 541 nsew
rlabel metal2 s 9546 10610 9654 10720 4 gnd
port 541 nsew
rlabel metal2 s 19530 4860 19638 4936 4 gnd
port 541 nsew
rlabel metal2 s 330 2174 438 2250 4 gnd
port 541 nsew
rlabel metal2 s 3306 21450 3414 21526 4 gnd
port 541 nsew
rlabel metal2 s 17034 23504 17142 23580 4 gnd
port 541 nsew
rlabel metal2 s 13290 19870 13398 19946 4 gnd
port 541 nsew
rlabel metal2 s 810 594 918 670 4 gnd
port 541 nsew
rlabel metal2 s 330 9820 438 9930 4 gnd
port 541 nsew
rlabel metal2 s 330 14560 438 14670 4 gnd
port 541 nsew
rlabel metal2 s 12042 15604 12150 15680 4 gnd
port 541 nsew
rlabel metal2 s 9546 1920 9654 2030 4 gnd
port 541 nsew
rlabel metal2 s 11562 10864 11670 10940 4 gnd
port 541 nsew
rlabel metal2 s 11562 14340 11670 14416 4 gnd
port 541 nsew
rlabel metal2 s 14058 21924 14166 22000 4 gnd
port 541 nsew
rlabel metal2 s 14538 16394 14646 16470 4 gnd
port 541 nsew
rlabel metal2 s 19050 3500 19158 3610 4 gnd
port 541 nsew
rlabel metal2 s 2058 11654 2166 11730 4 gnd
port 541 nsew
rlabel metal2 s 17802 24294 17910 24370 4 gnd
port 541 nsew
rlabel metal2 s 8298 2174 8406 2250 4 gnd
port 541 nsew
rlabel metal2 s 17034 15130 17142 15206 4 gnd
port 541 nsew
rlabel metal2 s 4074 12444 4182 12520 4 gnd
port 541 nsew
rlabel metal2 s 15306 17500 15414 17576 4 gnd
port 541 nsew
rlabel metal2 s 16554 18290 16662 18366 4 gnd
port 541 nsew
rlabel metal2 s 2058 10610 2166 10720 4 gnd
port 541 nsew
rlabel metal2 s 20298 1700 20406 1776 4 gnd
port 541 nsew
rlabel metal2 s 13290 19554 13398 19630 4 gnd
port 541 nsew
rlabel metal2 s 20298 16930 20406 17040 4 gnd
port 541 nsew
rlabel metal2 s 11562 7704 11670 7780 4 gnd
port 541 nsew
rlabel metal2 s 19530 18510 19638 18620 4 gnd
port 541 nsew
rlabel metal2 s 16554 17184 16662 17260 4 gnd
port 541 nsew
rlabel metal2 s 8298 17720 8406 17830 4 gnd
port 541 nsew
rlabel metal2 s 5322 1700 5430 1776 4 gnd
port 541 nsew
rlabel metal2 s 17802 1700 17910 1776 4 gnd
port 541 nsew
rlabel metal2 s 14058 3500 14166 3610 4 gnd
port 541 nsew
rlabel metal2 s 20298 10074 20406 10150 4 gnd
port 541 nsew
rlabel metal2 s 3306 23820 3414 23896 4 gnd
port 541 nsew
rlabel metal2 s 16554 19300 16662 19410 4 gnd
port 541 nsew
rlabel metal2 s 3306 2490 3414 2566 4 gnd
port 541 nsew
rlabel metal2 s 14058 10864 14166 10940 4 gnd
port 541 nsew
rlabel metal2 s 1578 13770 1686 13880 4 gnd
port 541 nsew
rlabel metal2 s 7818 16710 7926 16786 4 gnd
port 541 nsew
rlabel metal2 s 15306 25874 15414 25950 4 gnd
port 541 nsew
rlabel metal2 s 12810 3500 12918 3610 4 gnd
port 541 nsew
rlabel metal2 s 330 13550 438 13626 4 gnd
port 541 nsew
rlabel metal2 s 810 1384 918 1460 4 gnd
port 541 nsew
rlabel metal2 s 4554 8494 4662 8570 4 gnd
port 541 nsew
rlabel metal2 s 330 17720 438 17830 4 gnd
port 541 nsew
rlabel metal2 s 9066 2964 9174 3040 4 gnd
port 541 nsew
rlabel metal2 s 9066 14340 9174 14416 4 gnd
port 541 nsew
rlabel metal2 s 7050 25874 7158 25950 4 gnd
port 541 nsew
rlabel metal2 s 14538 21670 14646 21780 4 gnd
port 541 nsew
rlabel metal2 s 13290 4070 13398 4146 4 gnd
port 541 nsew
rlabel metal2 s 330 11654 438 11730 4 gnd
port 541 nsew
rlabel metal2 s 10794 10610 10902 10720 4 gnd
port 541 nsew
rlabel metal2 s 12810 19080 12918 19156 4 gnd
port 541 nsew
rlabel metal2 s 1578 20344 1686 20420 4 gnd
port 541 nsew
rlabel metal2 s 20778 9030 20886 9140 4 gnd
port 541 nsew
rlabel metal2 s 20778 3280 20886 3356 4 gnd
port 541 nsew
rlabel metal2 s 7050 12980 7158 13090 4 gnd
port 541 nsew
rlabel metal2 s 10314 15130 10422 15206 4 gnd
port 541 nsew
rlabel metal2 s 2826 2710 2934 2820 4 gnd
port 541 nsew
rlabel metal2 s 13290 16710 13398 16786 4 gnd
port 541 nsew
rlabel metal2 s 10794 11970 10902 12046 4 gnd
port 541 nsew
rlabel metal2 s 19530 8810 19638 8886 4 gnd
port 541 nsew
rlabel metal2 s 1578 18764 1686 18840 4 gnd
port 541 nsew
rlabel metal2 s 5322 23504 5430 23580 4 gnd
port 541 nsew
rlabel metal2 s 14058 8240 14166 8350 4 gnd
port 541 nsew
rlabel metal2 s 330 910 438 986 4 gnd
port 541 nsew
rlabel metal2 s 18282 19080 18390 19156 4 gnd
port 541 nsew
rlabel metal2 s 15786 11180 15894 11256 4 gnd
port 541 nsew
rlabel metal2 s 11562 2490 11670 2566 4 gnd
port 541 nsew
rlabel metal2 s 14538 19080 14646 19156 4 gnd
port 541 nsew
rlabel metal2 s 13290 1700 13398 1776 4 gnd
port 541 nsew
rlabel metal2 s 330 2710 438 2820 4 gnd
port 541 nsew
rlabel metal2 s 19050 14560 19158 14670 4 gnd
port 541 nsew
rlabel metal2 s 10794 14340 10902 14416 4 gnd
port 541 nsew
rlabel metal2 s 810 19870 918 19946 4 gnd
port 541 nsew
rlabel metal2 s 12810 15130 12918 15206 4 gnd
port 541 nsew
rlabel metal2 s 19050 1384 19158 1460 4 gnd
port 541 nsew
rlabel metal2 s 10314 1384 10422 1460 4 gnd
port 541 nsew
rlabel metal2 s 6570 25084 6678 25160 4 gnd
port 541 nsew
rlabel metal2 s 7818 11180 7926 11256 4 gnd
port 541 nsew
rlabel metal2 s 4554 21134 4662 21210 4 gnd
port 541 nsew
rlabel metal2 s 330 4070 438 4146 4 gnd
port 541 nsew
rlabel metal2 s 20778 20660 20886 20736 4 gnd
port 541 nsew
rlabel metal2 s 14538 4070 14646 4146 4 gnd
port 541 nsew
rlabel metal2 s 5802 14560 5910 14670 4 gnd
port 541 nsew
rlabel metal2 s 7818 2490 7926 2566 4 gnd
port 541 nsew
rlabel metal2 s 5802 8494 5910 8570 4 gnd
port 541 nsew
rlabel metal2 s 9066 24610 9174 24686 4 gnd
port 541 nsew
rlabel metal2 s 1578 9820 1686 9930 4 gnd
port 541 nsew
rlabel metal2 s 5322 7230 5430 7306 4 gnd
port 541 nsew
rlabel metal2 s 14058 8020 14166 8096 4 gnd
port 541 nsew
rlabel metal2 s 810 13550 918 13626 4 gnd
port 541 nsew
rlabel metal2 s 19050 1920 19158 2030 4 gnd
port 541 nsew
rlabel metal2 s 2058 25084 2166 25160 4 gnd
port 541 nsew
rlabel metal2 s 13290 15604 13398 15680 4 gnd
port 541 nsew
rlabel metal2 s 16554 20880 16662 20990 4 gnd
port 541 nsew
rlabel metal2 s 17802 13550 17910 13626 4 gnd
port 541 nsew
rlabel metal2 s 17802 5080 17910 5190 4 gnd
port 541 nsew
rlabel metal2 s 11562 8810 11670 8886 4 gnd
port 541 nsew
rlabel metal2 s 11562 12444 11670 12520 4 gnd
port 541 nsew
rlabel metal2 s 10314 4290 10422 4400 4 gnd
port 541 nsew
rlabel metal2 s 18282 11970 18390 12046 4 gnd
port 541 nsew
rlabel metal2 s 4074 23504 4182 23580 4 gnd
port 541 nsew
rlabel metal2 s 13290 8810 13398 8886 4 gnd
port 541 nsew
rlabel metal2 s 2826 4290 2934 4400 4 gnd
port 541 nsew
rlabel metal2 s 13290 16140 13398 16250 4 gnd
port 541 nsew
rlabel metal2 s 810 11970 918 12046 4 gnd
port 541 nsew
rlabel metal2 s 10794 1384 10902 1460 4 gnd
port 541 nsew
rlabel metal2 s 7818 6914 7926 6990 4 gnd
port 541 nsew
rlabel metal2 s 2826 23820 2934 23896 4 gnd
port 541 nsew
rlabel metal2 s 5322 21924 5430 22000 4 gnd
port 541 nsew
rlabel metal2 s 14538 17974 14646 18050 4 gnd
port 541 nsew
rlabel metal2 s 20298 20660 20406 20736 4 gnd
port 541 nsew
<< properties >>
string FIXED_BBOX 0 0 21216 26070
<< end >>
