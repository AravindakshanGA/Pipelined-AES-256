magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 2204 2731
<< nwell >>
rect -36 679 944 1471
<< pwell >>
rect 28 159 770 477
rect 28 25 874 159
<< scnmos >>
rect 114 51 144 451
rect 222 51 252 451
rect 330 51 360 451
rect 438 51 468 451
rect 546 51 576 451
rect 654 51 684 451
<< scpmos >>
rect 114 963 144 1363
rect 222 963 252 1363
rect 330 963 360 1363
rect 438 963 468 1363
rect 546 963 576 1363
rect 654 963 684 1363
<< ndiff >>
rect 54 268 114 451
rect 54 234 62 268
rect 96 234 114 268
rect 54 51 114 234
rect 144 268 222 451
rect 144 234 166 268
rect 200 234 222 268
rect 144 51 222 234
rect 252 268 330 451
rect 252 234 274 268
rect 308 234 330 268
rect 252 51 330 234
rect 360 268 438 451
rect 360 234 382 268
rect 416 234 438 268
rect 360 51 438 234
rect 468 268 546 451
rect 468 234 490 268
rect 524 234 546 268
rect 468 51 546 234
rect 576 268 654 451
rect 576 234 598 268
rect 632 234 654 268
rect 576 51 654 234
rect 684 268 744 451
rect 684 234 702 268
rect 736 234 744 268
rect 684 51 744 234
<< pdiff >>
rect 54 1180 114 1363
rect 54 1146 62 1180
rect 96 1146 114 1180
rect 54 963 114 1146
rect 144 1180 222 1363
rect 144 1146 166 1180
rect 200 1146 222 1180
rect 144 963 222 1146
rect 252 1180 330 1363
rect 252 1146 274 1180
rect 308 1146 330 1180
rect 252 963 330 1146
rect 360 1180 438 1363
rect 360 1146 382 1180
rect 416 1146 438 1180
rect 360 963 438 1146
rect 468 1180 546 1363
rect 468 1146 490 1180
rect 524 1146 546 1180
rect 468 963 546 1146
rect 576 1180 654 1363
rect 576 1146 598 1180
rect 632 1146 654 1180
rect 576 963 654 1146
rect 684 1180 744 1363
rect 684 1146 702 1180
rect 736 1146 744 1180
rect 684 963 744 1146
<< ndiffc >>
rect 62 234 96 268
rect 166 234 200 268
rect 274 234 308 268
rect 382 234 416 268
rect 490 234 524 268
rect 598 234 632 268
rect 702 234 736 268
<< pdiffc >>
rect 62 1146 96 1180
rect 166 1146 200 1180
rect 274 1146 308 1180
rect 382 1146 416 1180
rect 490 1146 524 1180
rect 598 1146 632 1180
rect 702 1146 736 1180
<< psubdiff >>
rect 798 109 848 133
rect 798 75 806 109
rect 840 75 848 109
rect 798 51 848 75
<< nsubdiff >>
rect 798 1326 848 1350
rect 798 1292 806 1326
rect 840 1292 848 1326
rect 798 1268 848 1292
<< psubdiffcont >>
rect 806 75 840 109
<< nsubdiffcont >>
rect 806 1292 840 1326
<< poly >>
rect 114 1363 144 1389
rect 222 1363 252 1389
rect 330 1363 360 1389
rect 438 1363 468 1389
rect 546 1363 576 1389
rect 654 1363 684 1389
rect 114 937 144 963
rect 222 937 252 963
rect 330 937 360 963
rect 438 937 468 963
rect 546 937 576 963
rect 654 937 684 963
rect 114 907 684 937
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
rect 114 477 684 507
rect 114 451 144 477
rect 222 451 252 477
rect 330 451 360 477
rect 438 451 468 477
rect 546 451 576 477
rect 654 451 684 477
rect 114 25 144 51
rect 222 25 252 51
rect 330 25 360 51
rect 438 25 468 51
rect 546 25 576 51
rect 654 25 684 51
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 908 1431
rect 62 1180 96 1397
rect 62 1130 96 1146
rect 166 1180 200 1196
rect 166 1096 200 1146
rect 274 1180 308 1397
rect 274 1130 308 1146
rect 382 1180 416 1196
rect 382 1096 416 1146
rect 490 1180 524 1397
rect 490 1130 524 1146
rect 598 1180 632 1196
rect 598 1096 632 1146
rect 702 1180 736 1397
rect 806 1326 840 1397
rect 806 1276 840 1292
rect 702 1130 736 1146
rect 166 1062 632 1096
rect 64 724 98 740
rect 64 674 98 690
rect 382 724 416 1062
rect 382 690 433 724
rect 382 352 416 690
rect 166 318 632 352
rect 62 268 96 284
rect 62 17 96 234
rect 166 268 200 318
rect 166 218 200 234
rect 274 268 308 284
rect 274 17 308 234
rect 382 268 416 318
rect 382 218 416 234
rect 490 268 524 284
rect 490 17 524 234
rect 598 268 632 318
rect 598 218 632 234
rect 702 268 736 284
rect 702 17 736 234
rect 806 109 840 125
rect 806 17 840 75
rect 0 -17 908 17
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 416 707 416 707 4 Z
port 2 nsew
rlabel locali s 454 0 454 0 4 gnd
port 3 nsew
rlabel locali s 454 1414 454 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 908 1079
<< end >>
