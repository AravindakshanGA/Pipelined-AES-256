magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1260 -1260 1261 1261
<< end >>
