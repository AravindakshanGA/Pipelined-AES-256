magic
tech sky130A
magscale 1 2
timestamp 1543373562
<< checkpaint >>
rect -1260 -1260 25066 28170
<< metal1 >>
rect 1517 0 1553 26910
rect 1589 0 1625 26910
rect 1733 0 1769 26910
rect 1805 0 1841 26910
rect 1997 0 2033 26910
rect 2069 0 2105 26910
rect 2213 0 2249 26910
rect 2285 0 2321 26910
rect 2765 0 2801 26910
rect 2837 0 2873 26910
rect 2981 0 3017 26910
rect 3053 0 3089 26910
rect 3245 0 3281 26910
rect 3317 0 3353 26910
rect 3461 0 3497 26910
rect 3533 0 3569 26910
rect 4013 0 4049 26910
rect 4085 0 4121 26910
rect 4229 0 4265 26910
rect 4301 0 4337 26910
rect 4493 0 4529 26910
rect 4565 0 4601 26910
rect 4709 0 4745 26910
rect 4781 0 4817 26910
rect 5261 0 5297 26910
rect 5333 0 5369 26910
rect 5477 0 5513 26910
rect 5549 0 5585 26910
rect 5741 0 5777 26910
rect 5813 0 5849 26910
rect 5957 0 5993 26910
rect 6029 0 6065 26910
rect 6509 0 6545 26910
rect 6581 0 6617 26910
rect 6725 0 6761 26910
rect 6797 0 6833 26910
rect 6989 0 7025 26910
rect 7061 0 7097 26910
rect 7205 0 7241 26910
rect 7277 0 7313 26910
rect 7757 0 7793 26910
rect 7829 0 7865 26910
rect 7973 0 8009 26910
rect 8045 0 8081 26910
rect 8237 0 8273 26910
rect 8309 0 8345 26910
rect 8453 0 8489 26910
rect 8525 0 8561 26910
rect 9005 0 9041 26910
rect 9077 0 9113 26910
rect 9221 0 9257 26910
rect 9293 0 9329 26910
rect 9485 0 9521 26910
rect 9557 0 9593 26910
rect 9701 0 9737 26910
rect 9773 0 9809 26910
rect 10253 0 10289 26910
rect 10325 0 10361 26910
rect 10469 0 10505 26910
rect 10541 0 10577 26910
rect 10733 0 10769 26910
rect 10805 0 10841 26910
rect 10949 0 10985 26910
rect 11021 0 11057 26910
rect 11501 0 11537 26910
rect 11573 0 11609 26910
rect 11717 0 11753 26910
rect 11789 0 11825 26910
rect 11981 0 12017 26910
rect 12053 0 12089 26910
rect 12197 0 12233 26910
rect 12269 0 12305 26910
rect 12749 0 12785 26910
rect 12821 0 12857 26910
rect 12965 0 13001 26910
rect 13037 0 13073 26910
rect 13229 0 13265 26910
rect 13301 0 13337 26910
rect 13445 0 13481 26910
rect 13517 0 13553 26910
rect 13997 0 14033 26910
rect 14069 0 14105 26910
rect 14213 0 14249 26910
rect 14285 0 14321 26910
rect 14477 0 14513 26910
rect 14549 0 14585 26910
rect 14693 0 14729 26910
rect 14765 0 14801 26910
rect 15245 0 15281 26910
rect 15317 0 15353 26910
rect 15461 0 15497 26910
rect 15533 0 15569 26910
rect 15725 0 15761 26910
rect 15797 0 15833 26910
rect 15941 0 15977 26910
rect 16013 0 16049 26910
rect 16493 0 16529 26910
rect 16565 0 16601 26910
rect 16709 0 16745 26910
rect 16781 0 16817 26910
rect 16973 0 17009 26910
rect 17045 0 17081 26910
rect 17189 0 17225 26910
rect 17261 0 17297 26910
rect 17741 0 17777 26910
rect 17813 0 17849 26910
rect 17957 0 17993 26910
rect 18029 0 18065 26910
rect 18221 0 18257 26910
rect 18293 0 18329 26910
rect 18437 0 18473 26910
rect 18509 0 18545 26910
rect 18989 0 19025 26910
rect 19061 0 19097 26910
rect 19205 0 19241 26910
rect 19277 0 19313 26910
rect 19469 0 19505 26910
rect 19541 0 19577 26910
rect 19685 0 19721 26910
rect 19757 0 19793 26910
rect 20237 0 20273 26910
rect 20309 0 20345 26910
rect 20453 0 20489 26910
rect 20525 0 20561 26910
rect 20717 0 20753 26910
rect 20789 0 20825 26910
rect 20933 0 20969 26910
rect 21005 0 21041 26910
rect 21485 0 21521 26910
rect 21557 0 21593 26910
rect 21701 0 21737 26910
rect 21773 0 21809 26910
rect 21965 0 22001 26910
rect 22037 0 22073 26910
rect 22181 0 22217 26910
rect 22253 0 22289 26910
<< metal2 >>
rect 38 26653 47 26709
rect 103 26695 112 26709
rect 23694 26695 23703 26709
rect 103 26667 23703 26695
rect 103 26653 112 26667
rect 23694 26653 23703 26667
rect 23759 26653 23768 26709
rect 448 26439 457 26495
rect 513 26481 522 26495
rect 23284 26481 23293 26495
rect 513 26453 23293 26481
rect 513 26439 522 26453
rect 23284 26439 23293 26453
rect 23349 26439 23358 26495
rect 621 26223 23185 26271
rect 448 26092 457 26148
rect 513 26134 522 26148
rect 23284 26134 23293 26148
rect 513 26106 23293 26134
rect 513 26092 522 26106
rect 23284 26092 23293 26106
rect 23349 26092 23358 26148
rect 621 25969 23185 26017
rect 448 25855 457 25911
rect 513 25897 522 25911
rect 23284 25897 23293 25911
rect 513 25869 23293 25897
rect 513 25855 522 25869
rect 23284 25855 23293 25869
rect 23349 25855 23358 25911
rect 621 25749 23185 25797
rect 621 25653 23185 25701
rect 448 25539 457 25595
rect 513 25581 522 25595
rect 23284 25581 23293 25595
rect 513 25553 23293 25581
rect 513 25539 522 25553
rect 23284 25539 23293 25553
rect 23349 25539 23358 25595
rect 621 25433 23185 25481
rect 448 25302 457 25358
rect 513 25344 522 25358
rect 23284 25344 23293 25358
rect 513 25316 23293 25344
rect 513 25302 522 25316
rect 23284 25302 23293 25316
rect 23349 25302 23358 25358
rect 621 25179 23185 25227
rect 448 25065 457 25121
rect 513 25107 522 25121
rect 23284 25107 23293 25121
rect 513 25079 23293 25107
rect 513 25065 522 25079
rect 23284 25065 23293 25079
rect 23349 25065 23358 25121
rect 621 24959 23185 25007
rect 621 24863 23185 24911
rect 448 24749 457 24805
rect 513 24791 522 24805
rect 23284 24791 23293 24805
rect 513 24763 23293 24791
rect 513 24749 522 24763
rect 23284 24749 23293 24763
rect 23349 24749 23358 24805
rect 621 24643 23185 24691
rect 448 24512 457 24568
rect 513 24554 522 24568
rect 23284 24554 23293 24568
rect 513 24526 23293 24554
rect 513 24512 522 24526
rect 23284 24512 23293 24526
rect 23349 24512 23358 24568
rect 621 24389 23185 24437
rect 448 24275 457 24331
rect 513 24317 522 24331
rect 23284 24317 23293 24331
rect 513 24289 23293 24317
rect 513 24275 522 24289
rect 23284 24275 23293 24289
rect 23349 24275 23358 24331
rect 621 24169 23185 24217
rect 621 24073 23185 24121
rect 448 23959 457 24015
rect 513 24001 522 24015
rect 23284 24001 23293 24015
rect 513 23973 23293 24001
rect 513 23959 522 23973
rect 23284 23959 23293 23973
rect 23349 23959 23358 24015
rect 621 23853 23185 23901
rect 448 23722 457 23778
rect 513 23764 522 23778
rect 23284 23764 23293 23778
rect 513 23736 23293 23764
rect 513 23722 522 23736
rect 23284 23722 23293 23736
rect 23349 23722 23358 23778
rect 621 23599 23185 23647
rect 448 23485 457 23541
rect 513 23527 522 23541
rect 23284 23527 23293 23541
rect 513 23499 23293 23527
rect 513 23485 522 23499
rect 23284 23485 23293 23499
rect 23349 23485 23358 23541
rect 621 23379 23185 23427
rect 621 23283 23185 23331
rect 448 23169 457 23225
rect 513 23211 522 23225
rect 23284 23211 23293 23225
rect 513 23183 23293 23211
rect 513 23169 522 23183
rect 23284 23169 23293 23183
rect 23349 23169 23358 23225
rect 621 23063 23185 23111
rect 448 22932 457 22988
rect 513 22974 522 22988
rect 23284 22974 23293 22988
rect 513 22946 23293 22974
rect 513 22932 522 22946
rect 23284 22932 23293 22946
rect 23349 22932 23358 22988
rect 621 22809 23185 22857
rect 448 22695 457 22751
rect 513 22737 522 22751
rect 23284 22737 23293 22751
rect 513 22709 23293 22737
rect 513 22695 522 22709
rect 23284 22695 23293 22709
rect 23349 22695 23358 22751
rect 621 22589 23185 22637
rect 621 22493 23185 22541
rect 448 22379 457 22435
rect 513 22421 522 22435
rect 23284 22421 23293 22435
rect 513 22393 23293 22421
rect 513 22379 522 22393
rect 23284 22379 23293 22393
rect 23349 22379 23358 22435
rect 621 22273 23185 22321
rect 448 22142 457 22198
rect 513 22184 522 22198
rect 23284 22184 23293 22198
rect 513 22156 23293 22184
rect 513 22142 522 22156
rect 23284 22142 23293 22156
rect 23349 22142 23358 22198
rect 621 22019 23185 22067
rect 448 21905 457 21961
rect 513 21947 522 21961
rect 23284 21947 23293 21961
rect 513 21919 23293 21947
rect 513 21905 522 21919
rect 23284 21905 23293 21919
rect 23349 21905 23358 21961
rect 621 21799 23185 21847
rect 621 21703 23185 21751
rect 448 21589 457 21645
rect 513 21631 522 21645
rect 23284 21631 23293 21645
rect 513 21603 23293 21631
rect 513 21589 522 21603
rect 23284 21589 23293 21603
rect 23349 21589 23358 21645
rect 621 21483 23185 21531
rect 448 21352 457 21408
rect 513 21394 522 21408
rect 23284 21394 23293 21408
rect 513 21366 23293 21394
rect 513 21352 522 21366
rect 23284 21352 23293 21366
rect 23349 21352 23358 21408
rect 621 21229 23185 21277
rect 448 21115 457 21171
rect 513 21157 522 21171
rect 23284 21157 23293 21171
rect 513 21129 23293 21157
rect 513 21115 522 21129
rect 23284 21115 23293 21129
rect 23349 21115 23358 21171
rect 621 21009 23185 21057
rect 621 20913 23185 20961
rect 448 20799 457 20855
rect 513 20841 522 20855
rect 23284 20841 23293 20855
rect 513 20813 23293 20841
rect 513 20799 522 20813
rect 23284 20799 23293 20813
rect 23349 20799 23358 20855
rect 621 20693 23185 20741
rect 448 20562 457 20618
rect 513 20604 522 20618
rect 23284 20604 23293 20618
rect 513 20576 23293 20604
rect 513 20562 522 20576
rect 23284 20562 23293 20576
rect 23349 20562 23358 20618
rect 621 20439 23185 20487
rect 448 20325 457 20381
rect 513 20367 522 20381
rect 23284 20367 23293 20381
rect 513 20339 23293 20367
rect 513 20325 522 20339
rect 23284 20325 23293 20339
rect 23349 20325 23358 20381
rect 621 20219 23185 20267
rect 621 20123 23185 20171
rect 448 20009 457 20065
rect 513 20051 522 20065
rect 23284 20051 23293 20065
rect 513 20023 23293 20051
rect 513 20009 522 20023
rect 23284 20009 23293 20023
rect 23349 20009 23358 20065
rect 621 19903 23185 19951
rect 448 19772 457 19828
rect 513 19814 522 19828
rect 23284 19814 23293 19828
rect 513 19786 23293 19814
rect 513 19772 522 19786
rect 23284 19772 23293 19786
rect 23349 19772 23358 19828
rect 621 19649 23185 19697
rect 448 19535 457 19591
rect 513 19577 522 19591
rect 23284 19577 23293 19591
rect 513 19549 23293 19577
rect 513 19535 522 19549
rect 23284 19535 23293 19549
rect 23349 19535 23358 19591
rect 621 19429 23185 19477
rect 621 19333 23185 19381
rect 448 19219 457 19275
rect 513 19261 522 19275
rect 23284 19261 23293 19275
rect 513 19233 23293 19261
rect 513 19219 522 19233
rect 23284 19219 23293 19233
rect 23349 19219 23358 19275
rect 621 19113 23185 19161
rect 448 18982 457 19038
rect 513 19024 522 19038
rect 23284 19024 23293 19038
rect 513 18996 23293 19024
rect 513 18982 522 18996
rect 23284 18982 23293 18996
rect 23349 18982 23358 19038
rect 621 18859 23185 18907
rect 448 18745 457 18801
rect 513 18787 522 18801
rect 23284 18787 23293 18801
rect 513 18759 23293 18787
rect 513 18745 522 18759
rect 23284 18745 23293 18759
rect 23349 18745 23358 18801
rect 621 18639 23185 18687
rect 621 18543 23185 18591
rect 448 18429 457 18485
rect 513 18471 522 18485
rect 23284 18471 23293 18485
rect 513 18443 23293 18471
rect 513 18429 522 18443
rect 23284 18429 23293 18443
rect 23349 18429 23358 18485
rect 621 18323 23185 18371
rect 448 18192 457 18248
rect 513 18234 522 18248
rect 23284 18234 23293 18248
rect 513 18206 23293 18234
rect 513 18192 522 18206
rect 23284 18192 23293 18206
rect 23349 18192 23358 18248
rect 621 18069 23185 18117
rect 448 17955 457 18011
rect 513 17997 522 18011
rect 23284 17997 23293 18011
rect 513 17969 23293 17997
rect 513 17955 522 17969
rect 23284 17955 23293 17969
rect 23349 17955 23358 18011
rect 621 17849 23185 17897
rect 621 17753 23185 17801
rect 448 17639 457 17695
rect 513 17681 522 17695
rect 23284 17681 23293 17695
rect 513 17653 23293 17681
rect 513 17639 522 17653
rect 23284 17639 23293 17653
rect 23349 17639 23358 17695
rect 621 17533 23185 17581
rect 448 17402 457 17458
rect 513 17444 522 17458
rect 23284 17444 23293 17458
rect 513 17416 23293 17444
rect 513 17402 522 17416
rect 23284 17402 23293 17416
rect 23349 17402 23358 17458
rect 621 17279 23185 17327
rect 448 17165 457 17221
rect 513 17207 522 17221
rect 23284 17207 23293 17221
rect 513 17179 23293 17207
rect 513 17165 522 17179
rect 23284 17165 23293 17179
rect 23349 17165 23358 17221
rect 621 17059 23185 17107
rect 621 16963 23185 17011
rect 448 16849 457 16905
rect 513 16891 522 16905
rect 23284 16891 23293 16905
rect 513 16863 23293 16891
rect 513 16849 522 16863
rect 23284 16849 23293 16863
rect 23349 16849 23358 16905
rect 621 16743 23185 16791
rect 448 16612 457 16668
rect 513 16654 522 16668
rect 23284 16654 23293 16668
rect 513 16626 23293 16654
rect 513 16612 522 16626
rect 23284 16612 23293 16626
rect 23349 16612 23358 16668
rect 621 16489 23185 16537
rect 448 16375 457 16431
rect 513 16417 522 16431
rect 23284 16417 23293 16431
rect 513 16389 23293 16417
rect 513 16375 522 16389
rect 23284 16375 23293 16389
rect 23349 16375 23358 16431
rect 621 16269 23185 16317
rect 621 16173 23185 16221
rect 448 16059 457 16115
rect 513 16101 522 16115
rect 23284 16101 23293 16115
rect 513 16073 23293 16101
rect 513 16059 522 16073
rect 23284 16059 23293 16073
rect 23349 16059 23358 16115
rect 621 15953 23185 16001
rect 448 15822 457 15878
rect 513 15864 522 15878
rect 23284 15864 23293 15878
rect 513 15836 23293 15864
rect 513 15822 522 15836
rect 23284 15822 23293 15836
rect 23349 15822 23358 15878
rect 621 15699 23185 15747
rect 448 15585 457 15641
rect 513 15627 522 15641
rect 23284 15627 23293 15641
rect 513 15599 23293 15627
rect 513 15585 522 15599
rect 23284 15585 23293 15599
rect 23349 15585 23358 15641
rect 621 15479 23185 15527
rect 621 15383 23185 15431
rect 448 15269 457 15325
rect 513 15311 522 15325
rect 23284 15311 23293 15325
rect 513 15283 23293 15311
rect 513 15269 522 15283
rect 23284 15269 23293 15283
rect 23349 15269 23358 15325
rect 621 15163 23185 15211
rect 448 15032 457 15088
rect 513 15074 522 15088
rect 23284 15074 23293 15088
rect 513 15046 23293 15074
rect 513 15032 522 15046
rect 23284 15032 23293 15046
rect 23349 15032 23358 15088
rect 621 14909 23185 14957
rect 448 14795 457 14851
rect 513 14837 522 14851
rect 23284 14837 23293 14851
rect 513 14809 23293 14837
rect 513 14795 522 14809
rect 23284 14795 23293 14809
rect 23349 14795 23358 14851
rect 621 14689 23185 14737
rect 621 14593 23185 14641
rect 448 14479 457 14535
rect 513 14521 522 14535
rect 23284 14521 23293 14535
rect 513 14493 23293 14521
rect 513 14479 522 14493
rect 23284 14479 23293 14493
rect 23349 14479 23358 14535
rect 621 14373 23185 14421
rect 448 14242 457 14298
rect 513 14284 522 14298
rect 23284 14284 23293 14298
rect 513 14256 23293 14284
rect 513 14242 522 14256
rect 23284 14242 23293 14256
rect 23349 14242 23358 14298
rect 621 14119 23185 14167
rect 448 14005 457 14061
rect 513 14047 522 14061
rect 23284 14047 23293 14061
rect 513 14019 23293 14047
rect 513 14005 522 14019
rect 23284 14005 23293 14019
rect 23349 14005 23358 14061
rect 621 13899 23185 13947
rect 621 13803 23185 13851
rect 448 13689 457 13745
rect 513 13731 522 13745
rect 23284 13731 23293 13745
rect 513 13703 23293 13731
rect 513 13689 522 13703
rect 23284 13689 23293 13703
rect 23349 13689 23358 13745
rect 621 13583 23185 13631
rect 448 13452 457 13508
rect 513 13494 522 13508
rect 23284 13494 23293 13508
rect 513 13466 23293 13494
rect 513 13452 522 13466
rect 23284 13452 23293 13466
rect 23349 13452 23358 13508
rect 621 13329 23185 13377
rect 448 13215 457 13271
rect 513 13257 522 13271
rect 23284 13257 23293 13271
rect 513 13229 23293 13257
rect 513 13215 522 13229
rect 23284 13215 23293 13229
rect 23349 13215 23358 13271
rect 621 13109 23185 13157
rect 621 13013 23185 13061
rect 448 12899 457 12955
rect 513 12941 522 12955
rect 23284 12941 23293 12955
rect 513 12913 23293 12941
rect 513 12899 522 12913
rect 23284 12899 23293 12913
rect 23349 12899 23358 12955
rect 621 12793 23185 12841
rect 448 12662 457 12718
rect 513 12704 522 12718
rect 23284 12704 23293 12718
rect 513 12676 23293 12704
rect 513 12662 522 12676
rect 23284 12662 23293 12676
rect 23349 12662 23358 12718
rect 621 12539 23185 12587
rect 448 12425 457 12481
rect 513 12467 522 12481
rect 23284 12467 23293 12481
rect 513 12439 23293 12467
rect 513 12425 522 12439
rect 23284 12425 23293 12439
rect 23349 12425 23358 12481
rect 621 12319 23185 12367
rect 621 12223 23185 12271
rect 448 12109 457 12165
rect 513 12151 522 12165
rect 23284 12151 23293 12165
rect 513 12123 23293 12151
rect 513 12109 522 12123
rect 23284 12109 23293 12123
rect 23349 12109 23358 12165
rect 621 12003 23185 12051
rect 448 11872 457 11928
rect 513 11914 522 11928
rect 23284 11914 23293 11928
rect 513 11886 23293 11914
rect 513 11872 522 11886
rect 23284 11872 23293 11886
rect 23349 11872 23358 11928
rect 621 11749 23185 11797
rect 448 11635 457 11691
rect 513 11677 522 11691
rect 23284 11677 23293 11691
rect 513 11649 23293 11677
rect 513 11635 522 11649
rect 23284 11635 23293 11649
rect 23349 11635 23358 11691
rect 621 11529 23185 11577
rect 621 11433 23185 11481
rect 448 11319 457 11375
rect 513 11361 522 11375
rect 23284 11361 23293 11375
rect 513 11333 23293 11361
rect 513 11319 522 11333
rect 23284 11319 23293 11333
rect 23349 11319 23358 11375
rect 621 11213 23185 11261
rect 448 11082 457 11138
rect 513 11124 522 11138
rect 23284 11124 23293 11138
rect 513 11096 23293 11124
rect 513 11082 522 11096
rect 23284 11082 23293 11096
rect 23349 11082 23358 11138
rect 621 10959 23185 11007
rect 448 10845 457 10901
rect 513 10887 522 10901
rect 23284 10887 23293 10901
rect 513 10859 23293 10887
rect 513 10845 522 10859
rect 23284 10845 23293 10859
rect 23349 10845 23358 10901
rect 621 10739 23185 10787
rect 621 10643 23185 10691
rect 448 10529 457 10585
rect 513 10571 522 10585
rect 23284 10571 23293 10585
rect 513 10543 23293 10571
rect 513 10529 522 10543
rect 23284 10529 23293 10543
rect 23349 10529 23358 10585
rect 621 10423 23185 10471
rect 448 10292 457 10348
rect 513 10334 522 10348
rect 23284 10334 23293 10348
rect 513 10306 23293 10334
rect 513 10292 522 10306
rect 23284 10292 23293 10306
rect 23349 10292 23358 10348
rect 621 10169 23185 10217
rect 448 10055 457 10111
rect 513 10097 522 10111
rect 23284 10097 23293 10111
rect 513 10069 23293 10097
rect 513 10055 522 10069
rect 23284 10055 23293 10069
rect 23349 10055 23358 10111
rect 621 9949 23185 9997
rect 621 9853 23185 9901
rect 448 9739 457 9795
rect 513 9781 522 9795
rect 23284 9781 23293 9795
rect 513 9753 23293 9781
rect 513 9739 522 9753
rect 23284 9739 23293 9753
rect 23349 9739 23358 9795
rect 621 9633 23185 9681
rect 448 9502 457 9558
rect 513 9544 522 9558
rect 23284 9544 23293 9558
rect 513 9516 23293 9544
rect 513 9502 522 9516
rect 23284 9502 23293 9516
rect 23349 9502 23358 9558
rect 621 9379 23185 9427
rect 448 9265 457 9321
rect 513 9307 522 9321
rect 23284 9307 23293 9321
rect 513 9279 23293 9307
rect 513 9265 522 9279
rect 23284 9265 23293 9279
rect 23349 9265 23358 9321
rect 621 9159 23185 9207
rect 621 9063 23185 9111
rect 448 8949 457 9005
rect 513 8991 522 9005
rect 23284 8991 23293 9005
rect 513 8963 23293 8991
rect 513 8949 522 8963
rect 23284 8949 23293 8963
rect 23349 8949 23358 9005
rect 621 8843 23185 8891
rect 448 8712 457 8768
rect 513 8754 522 8768
rect 23284 8754 23293 8768
rect 513 8726 23293 8754
rect 513 8712 522 8726
rect 23284 8712 23293 8726
rect 23349 8712 23358 8768
rect 621 8589 23185 8637
rect 448 8475 457 8531
rect 513 8517 522 8531
rect 23284 8517 23293 8531
rect 513 8489 23293 8517
rect 513 8475 522 8489
rect 23284 8475 23293 8489
rect 23349 8475 23358 8531
rect 621 8369 23185 8417
rect 621 8273 23185 8321
rect 448 8159 457 8215
rect 513 8201 522 8215
rect 23284 8201 23293 8215
rect 513 8173 23293 8201
rect 513 8159 522 8173
rect 23284 8159 23293 8173
rect 23349 8159 23358 8215
rect 621 8053 23185 8101
rect 448 7922 457 7978
rect 513 7964 522 7978
rect 23284 7964 23293 7978
rect 513 7936 23293 7964
rect 513 7922 522 7936
rect 23284 7922 23293 7936
rect 23349 7922 23358 7978
rect 621 7799 23185 7847
rect 448 7685 457 7741
rect 513 7727 522 7741
rect 23284 7727 23293 7741
rect 513 7699 23293 7727
rect 513 7685 522 7699
rect 23284 7685 23293 7699
rect 23349 7685 23358 7741
rect 621 7579 23185 7627
rect 621 7483 23185 7531
rect 448 7369 457 7425
rect 513 7411 522 7425
rect 23284 7411 23293 7425
rect 513 7383 23293 7411
rect 513 7369 522 7383
rect 23284 7369 23293 7383
rect 23349 7369 23358 7425
rect 621 7263 23185 7311
rect 448 7132 457 7188
rect 513 7174 522 7188
rect 23284 7174 23293 7188
rect 513 7146 23293 7174
rect 513 7132 522 7146
rect 23284 7132 23293 7146
rect 23349 7132 23358 7188
rect 621 7009 23185 7057
rect 448 6895 457 6951
rect 513 6937 522 6951
rect 23284 6937 23293 6951
rect 513 6909 23293 6937
rect 513 6895 522 6909
rect 23284 6895 23293 6909
rect 23349 6895 23358 6951
rect 621 6789 23185 6837
rect 621 6693 23185 6741
rect 448 6579 457 6635
rect 513 6621 522 6635
rect 23284 6621 23293 6635
rect 513 6593 23293 6621
rect 513 6579 522 6593
rect 23284 6579 23293 6593
rect 23349 6579 23358 6635
rect 621 6473 23185 6521
rect 448 6342 457 6398
rect 513 6384 522 6398
rect 23284 6384 23293 6398
rect 513 6356 23293 6384
rect 513 6342 522 6356
rect 23284 6342 23293 6356
rect 23349 6342 23358 6398
rect 621 6219 23185 6267
rect 448 6105 457 6161
rect 513 6147 522 6161
rect 23284 6147 23293 6161
rect 513 6119 23293 6147
rect 513 6105 522 6119
rect 23284 6105 23293 6119
rect 23349 6105 23358 6161
rect 621 5999 23185 6047
rect 621 5903 23185 5951
rect 448 5789 457 5845
rect 513 5831 522 5845
rect 23284 5831 23293 5845
rect 513 5803 23293 5831
rect 513 5789 522 5803
rect 23284 5789 23293 5803
rect 23349 5789 23358 5845
rect 621 5683 23185 5731
rect 448 5552 457 5608
rect 513 5594 522 5608
rect 23284 5594 23293 5608
rect 513 5566 23293 5594
rect 513 5552 522 5566
rect 23284 5552 23293 5566
rect 23349 5552 23358 5608
rect 621 5429 23185 5477
rect 448 5315 457 5371
rect 513 5357 522 5371
rect 23284 5357 23293 5371
rect 513 5329 23293 5357
rect 513 5315 522 5329
rect 23284 5315 23293 5329
rect 23349 5315 23358 5371
rect 621 5209 23185 5257
rect 621 5113 23185 5161
rect 448 4999 457 5055
rect 513 5041 522 5055
rect 23284 5041 23293 5055
rect 513 5013 23293 5041
rect 513 4999 522 5013
rect 23284 4999 23293 5013
rect 23349 4999 23358 5055
rect 621 4893 23185 4941
rect 448 4762 457 4818
rect 513 4804 522 4818
rect 23284 4804 23293 4818
rect 513 4776 23293 4804
rect 513 4762 522 4776
rect 23284 4762 23293 4776
rect 23349 4762 23358 4818
rect 621 4639 23185 4687
rect 448 4525 457 4581
rect 513 4567 522 4581
rect 23284 4567 23293 4581
rect 513 4539 23293 4567
rect 513 4525 522 4539
rect 23284 4525 23293 4539
rect 23349 4525 23358 4581
rect 621 4419 23185 4467
rect 621 4323 23185 4371
rect 448 4209 457 4265
rect 513 4251 522 4265
rect 23284 4251 23293 4265
rect 513 4223 23293 4251
rect 513 4209 522 4223
rect 23284 4209 23293 4223
rect 23349 4209 23358 4265
rect 621 4103 23185 4151
rect 448 3972 457 4028
rect 513 4014 522 4028
rect 23284 4014 23293 4028
rect 513 3986 23293 4014
rect 513 3972 522 3986
rect 23284 3972 23293 3986
rect 23349 3972 23358 4028
rect 621 3849 23185 3897
rect 448 3735 457 3791
rect 513 3777 522 3791
rect 23284 3777 23293 3791
rect 513 3749 23293 3777
rect 513 3735 522 3749
rect 23284 3735 23293 3749
rect 23349 3735 23358 3791
rect 621 3629 23185 3677
rect 621 3533 23185 3581
rect 448 3419 457 3475
rect 513 3461 522 3475
rect 23284 3461 23293 3475
rect 513 3433 23293 3461
rect 513 3419 522 3433
rect 23284 3419 23293 3433
rect 23349 3419 23358 3475
rect 621 3313 23185 3361
rect 448 3182 457 3238
rect 513 3224 522 3238
rect 23284 3224 23293 3238
rect 513 3196 23293 3224
rect 513 3182 522 3196
rect 23284 3182 23293 3196
rect 23349 3182 23358 3238
rect 621 3059 23185 3107
rect 448 2945 457 3001
rect 513 2987 522 3001
rect 23284 2987 23293 3001
rect 513 2959 23293 2987
rect 513 2945 522 2959
rect 23284 2945 23293 2959
rect 23349 2945 23358 3001
rect 621 2839 23185 2887
rect 621 2743 23185 2791
rect 448 2629 457 2685
rect 513 2671 522 2685
rect 23284 2671 23293 2685
rect 513 2643 23293 2671
rect 513 2629 522 2643
rect 23284 2629 23293 2643
rect 23349 2629 23358 2685
rect 621 2523 23185 2571
rect 448 2392 457 2448
rect 513 2434 522 2448
rect 23284 2434 23293 2448
rect 513 2406 23293 2434
rect 513 2392 522 2406
rect 23284 2392 23293 2406
rect 23349 2392 23358 2448
rect 621 2269 23185 2317
rect 448 2155 457 2211
rect 513 2197 522 2211
rect 23284 2197 23293 2211
rect 513 2169 23293 2197
rect 513 2155 522 2169
rect 23284 2155 23293 2169
rect 23349 2155 23358 2211
rect 621 2049 23185 2097
rect 621 1953 23185 2001
rect 448 1839 457 1895
rect 513 1881 522 1895
rect 23284 1881 23293 1895
rect 513 1853 23293 1881
rect 513 1839 522 1853
rect 23284 1839 23293 1853
rect 23349 1839 23358 1895
rect 621 1733 23185 1781
rect 448 1602 457 1658
rect 513 1644 522 1658
rect 23284 1644 23293 1658
rect 513 1616 23293 1644
rect 513 1602 522 1616
rect 23284 1602 23293 1616
rect 23349 1602 23358 1658
rect 621 1479 23185 1527
rect 448 1365 457 1421
rect 513 1407 522 1421
rect 23284 1407 23293 1421
rect 513 1379 23293 1407
rect 513 1365 522 1379
rect 23284 1365 23293 1379
rect 23349 1365 23358 1421
rect 621 1259 23185 1307
rect 621 1163 23185 1211
rect 448 1049 457 1105
rect 513 1091 522 1105
rect 23284 1091 23293 1105
rect 513 1063 23293 1091
rect 513 1049 522 1063
rect 23284 1049 23293 1063
rect 23349 1049 23358 1105
rect 621 943 23185 991
rect 448 812 457 868
rect 513 854 522 868
rect 23284 854 23293 868
rect 513 826 23293 854
rect 513 812 522 826
rect 23284 812 23293 826
rect 23349 812 23358 868
rect 448 685 457 741
rect 513 727 522 741
rect 23284 727 23293 741
rect 513 699 23293 727
rect 513 685 522 699
rect 23284 685 23293 699
rect 23349 685 23358 741
rect 621 469 23185 517
rect 38 251 47 307
rect 103 293 112 307
rect 23694 293 23703 307
rect 103 265 23703 293
rect 103 251 112 265
rect 23694 251 23703 265
rect 23759 251 23768 307
<< via2 >>
rect 47 26653 103 26709
rect 23703 26653 23759 26709
rect 457 26439 513 26495
rect 23293 26439 23349 26495
rect 457 26092 513 26148
rect 23293 26092 23349 26148
rect 457 25855 513 25911
rect 23293 25855 23349 25911
rect 457 25539 513 25595
rect 23293 25539 23349 25595
rect 457 25302 513 25358
rect 23293 25302 23349 25358
rect 457 25065 513 25121
rect 23293 25065 23349 25121
rect 457 24749 513 24805
rect 23293 24749 23349 24805
rect 457 24512 513 24568
rect 23293 24512 23349 24568
rect 457 24275 513 24331
rect 23293 24275 23349 24331
rect 457 23959 513 24015
rect 23293 23959 23349 24015
rect 457 23722 513 23778
rect 23293 23722 23349 23778
rect 457 23485 513 23541
rect 23293 23485 23349 23541
rect 457 23169 513 23225
rect 23293 23169 23349 23225
rect 457 22932 513 22988
rect 23293 22932 23349 22988
rect 457 22695 513 22751
rect 23293 22695 23349 22751
rect 457 22379 513 22435
rect 23293 22379 23349 22435
rect 457 22142 513 22198
rect 23293 22142 23349 22198
rect 457 21905 513 21961
rect 23293 21905 23349 21961
rect 457 21589 513 21645
rect 23293 21589 23349 21645
rect 457 21352 513 21408
rect 23293 21352 23349 21408
rect 457 21115 513 21171
rect 23293 21115 23349 21171
rect 457 20799 513 20855
rect 23293 20799 23349 20855
rect 457 20562 513 20618
rect 23293 20562 23349 20618
rect 457 20325 513 20381
rect 23293 20325 23349 20381
rect 457 20009 513 20065
rect 23293 20009 23349 20065
rect 457 19772 513 19828
rect 23293 19772 23349 19828
rect 457 19535 513 19591
rect 23293 19535 23349 19591
rect 457 19219 513 19275
rect 23293 19219 23349 19275
rect 457 18982 513 19038
rect 23293 18982 23349 19038
rect 457 18745 513 18801
rect 23293 18745 23349 18801
rect 457 18429 513 18485
rect 23293 18429 23349 18485
rect 457 18192 513 18248
rect 23293 18192 23349 18248
rect 457 17955 513 18011
rect 23293 17955 23349 18011
rect 457 17639 513 17695
rect 23293 17639 23349 17695
rect 457 17402 513 17458
rect 23293 17402 23349 17458
rect 457 17165 513 17221
rect 23293 17165 23349 17221
rect 457 16849 513 16905
rect 23293 16849 23349 16905
rect 457 16612 513 16668
rect 23293 16612 23349 16668
rect 457 16375 513 16431
rect 23293 16375 23349 16431
rect 457 16059 513 16115
rect 23293 16059 23349 16115
rect 457 15822 513 15878
rect 23293 15822 23349 15878
rect 457 15585 513 15641
rect 23293 15585 23349 15641
rect 457 15269 513 15325
rect 23293 15269 23349 15325
rect 457 15032 513 15088
rect 23293 15032 23349 15088
rect 457 14795 513 14851
rect 23293 14795 23349 14851
rect 457 14479 513 14535
rect 23293 14479 23349 14535
rect 457 14242 513 14298
rect 23293 14242 23349 14298
rect 457 14005 513 14061
rect 23293 14005 23349 14061
rect 457 13689 513 13745
rect 23293 13689 23349 13745
rect 457 13452 513 13508
rect 23293 13452 23349 13508
rect 457 13215 513 13271
rect 23293 13215 23349 13271
rect 457 12899 513 12955
rect 23293 12899 23349 12955
rect 457 12662 513 12718
rect 23293 12662 23349 12718
rect 457 12425 513 12481
rect 23293 12425 23349 12481
rect 457 12109 513 12165
rect 23293 12109 23349 12165
rect 457 11872 513 11928
rect 23293 11872 23349 11928
rect 457 11635 513 11691
rect 23293 11635 23349 11691
rect 457 11319 513 11375
rect 23293 11319 23349 11375
rect 457 11082 513 11138
rect 23293 11082 23349 11138
rect 457 10845 513 10901
rect 23293 10845 23349 10901
rect 457 10529 513 10585
rect 23293 10529 23349 10585
rect 457 10292 513 10348
rect 23293 10292 23349 10348
rect 457 10055 513 10111
rect 23293 10055 23349 10111
rect 457 9739 513 9795
rect 23293 9739 23349 9795
rect 457 9502 513 9558
rect 23293 9502 23349 9558
rect 457 9265 513 9321
rect 23293 9265 23349 9321
rect 457 8949 513 9005
rect 23293 8949 23349 9005
rect 457 8712 513 8768
rect 23293 8712 23349 8768
rect 457 8475 513 8531
rect 23293 8475 23349 8531
rect 457 8159 513 8215
rect 23293 8159 23349 8215
rect 457 7922 513 7978
rect 23293 7922 23349 7978
rect 457 7685 513 7741
rect 23293 7685 23349 7741
rect 457 7369 513 7425
rect 23293 7369 23349 7425
rect 457 7132 513 7188
rect 23293 7132 23349 7188
rect 457 6895 513 6951
rect 23293 6895 23349 6951
rect 457 6579 513 6635
rect 23293 6579 23349 6635
rect 457 6342 513 6398
rect 23293 6342 23349 6398
rect 457 6105 513 6161
rect 23293 6105 23349 6161
rect 457 5789 513 5845
rect 23293 5789 23349 5845
rect 457 5552 513 5608
rect 23293 5552 23349 5608
rect 457 5315 513 5371
rect 23293 5315 23349 5371
rect 457 4999 513 5055
rect 23293 4999 23349 5055
rect 457 4762 513 4818
rect 23293 4762 23349 4818
rect 457 4525 513 4581
rect 23293 4525 23349 4581
rect 457 4209 513 4265
rect 23293 4209 23349 4265
rect 457 3972 513 4028
rect 23293 3972 23349 4028
rect 457 3735 513 3791
rect 23293 3735 23349 3791
rect 457 3419 513 3475
rect 23293 3419 23349 3475
rect 457 3182 513 3238
rect 23293 3182 23349 3238
rect 457 2945 513 3001
rect 23293 2945 23349 3001
rect 457 2629 513 2685
rect 23293 2629 23349 2685
rect 457 2392 513 2448
rect 23293 2392 23349 2448
rect 457 2155 513 2211
rect 23293 2155 23349 2211
rect 457 1839 513 1895
rect 23293 1839 23349 1895
rect 457 1602 513 1658
rect 23293 1602 23349 1658
rect 457 1365 513 1421
rect 23293 1365 23349 1421
rect 457 1049 513 1105
rect 23293 1049 23349 1105
rect 457 812 513 868
rect 23293 812 23349 868
rect 457 685 513 741
rect 23293 685 23349 741
rect 47 251 103 307
rect 23703 251 23759 307
<< metal3 >>
rect 42 26713 108 26714
rect 23698 26713 23764 26714
rect 0 26649 43 26713
rect 107 26649 150 26713
rect 23656 26649 23699 26713
rect 23763 26649 23806 26713
rect 42 26648 108 26649
rect 23698 26648 23764 26649
rect 452 26499 518 26500
rect 23288 26499 23354 26500
rect 410 26435 453 26499
rect 517 26435 560 26499
rect 23246 26435 23289 26499
rect 23353 26435 23396 26499
rect 452 26434 518 26435
rect 23288 26434 23354 26435
rect 452 26152 518 26153
rect 23288 26152 23354 26153
rect 410 26088 453 26152
rect 517 26088 560 26152
rect 23246 26088 23289 26152
rect 23353 26088 23396 26152
rect 452 26087 518 26088
rect 23288 26087 23354 26088
rect 452 25915 518 25916
rect 23288 25915 23354 25916
rect 410 25851 453 25915
rect 517 25851 560 25915
rect 23246 25851 23289 25915
rect 23353 25851 23396 25915
rect 452 25850 518 25851
rect 23288 25850 23354 25851
rect 452 25599 518 25600
rect 23288 25599 23354 25600
rect 410 25535 453 25599
rect 517 25535 560 25599
rect 23246 25535 23289 25599
rect 23353 25535 23396 25599
rect 452 25534 518 25535
rect 23288 25534 23354 25535
rect 452 25362 518 25363
rect 23288 25362 23354 25363
rect 410 25298 453 25362
rect 517 25298 560 25362
rect 23246 25298 23289 25362
rect 23353 25298 23396 25362
rect 452 25297 518 25298
rect 23288 25297 23354 25298
rect 452 25125 518 25126
rect 23288 25125 23354 25126
rect 410 25061 453 25125
rect 517 25061 560 25125
rect 23246 25061 23289 25125
rect 23353 25061 23396 25125
rect 452 25060 518 25061
rect 23288 25060 23354 25061
rect 452 24809 518 24810
rect 23288 24809 23354 24810
rect 410 24745 453 24809
rect 517 24745 560 24809
rect 23246 24745 23289 24809
rect 23353 24745 23396 24809
rect 452 24744 518 24745
rect 23288 24744 23354 24745
rect 452 24572 518 24573
rect 23288 24572 23354 24573
rect 410 24508 453 24572
rect 517 24508 560 24572
rect 23246 24508 23289 24572
rect 23353 24508 23396 24572
rect 452 24507 518 24508
rect 23288 24507 23354 24508
rect 452 24335 518 24336
rect 23288 24335 23354 24336
rect 410 24271 453 24335
rect 517 24271 560 24335
rect 23246 24271 23289 24335
rect 23353 24271 23396 24335
rect 452 24270 518 24271
rect 23288 24270 23354 24271
rect 452 24019 518 24020
rect 23288 24019 23354 24020
rect 410 23955 453 24019
rect 517 23955 560 24019
rect 23246 23955 23289 24019
rect 23353 23955 23396 24019
rect 452 23954 518 23955
rect 23288 23954 23354 23955
rect 452 23782 518 23783
rect 23288 23782 23354 23783
rect 410 23718 453 23782
rect 517 23718 560 23782
rect 23246 23718 23289 23782
rect 23353 23718 23396 23782
rect 452 23717 518 23718
rect 23288 23717 23354 23718
rect 452 23545 518 23546
rect 23288 23545 23354 23546
rect 410 23481 453 23545
rect 517 23481 560 23545
rect 23246 23481 23289 23545
rect 23353 23481 23396 23545
rect 452 23480 518 23481
rect 23288 23480 23354 23481
rect 452 23229 518 23230
rect 23288 23229 23354 23230
rect 410 23165 453 23229
rect 517 23165 560 23229
rect 23246 23165 23289 23229
rect 23353 23165 23396 23229
rect 452 23164 518 23165
rect 23288 23164 23354 23165
rect 452 22992 518 22993
rect 23288 22992 23354 22993
rect 410 22928 453 22992
rect 517 22928 560 22992
rect 23246 22928 23289 22992
rect 23353 22928 23396 22992
rect 452 22927 518 22928
rect 23288 22927 23354 22928
rect 452 22755 518 22756
rect 23288 22755 23354 22756
rect 410 22691 453 22755
rect 517 22691 560 22755
rect 23246 22691 23289 22755
rect 23353 22691 23396 22755
rect 452 22690 518 22691
rect 23288 22690 23354 22691
rect 452 22439 518 22440
rect 23288 22439 23354 22440
rect 410 22375 453 22439
rect 517 22375 560 22439
rect 23246 22375 23289 22439
rect 23353 22375 23396 22439
rect 452 22374 518 22375
rect 23288 22374 23354 22375
rect 452 22202 518 22203
rect 23288 22202 23354 22203
rect 410 22138 453 22202
rect 517 22138 560 22202
rect 23246 22138 23289 22202
rect 23353 22138 23396 22202
rect 452 22137 518 22138
rect 23288 22137 23354 22138
rect 452 21965 518 21966
rect 23288 21965 23354 21966
rect 410 21901 453 21965
rect 517 21901 560 21965
rect 23246 21901 23289 21965
rect 23353 21901 23396 21965
rect 452 21900 518 21901
rect 23288 21900 23354 21901
rect 452 21649 518 21650
rect 23288 21649 23354 21650
rect 410 21585 453 21649
rect 517 21585 560 21649
rect 23246 21585 23289 21649
rect 23353 21585 23396 21649
rect 452 21584 518 21585
rect 23288 21584 23354 21585
rect 452 21412 518 21413
rect 23288 21412 23354 21413
rect 410 21348 453 21412
rect 517 21348 560 21412
rect 23246 21348 23289 21412
rect 23353 21348 23396 21412
rect 452 21347 518 21348
rect 23288 21347 23354 21348
rect 452 21175 518 21176
rect 23288 21175 23354 21176
rect 410 21111 453 21175
rect 517 21111 560 21175
rect 23246 21111 23289 21175
rect 23353 21111 23396 21175
rect 452 21110 518 21111
rect 23288 21110 23354 21111
rect 452 20859 518 20860
rect 23288 20859 23354 20860
rect 410 20795 453 20859
rect 517 20795 560 20859
rect 23246 20795 23289 20859
rect 23353 20795 23396 20859
rect 452 20794 518 20795
rect 23288 20794 23354 20795
rect 452 20622 518 20623
rect 23288 20622 23354 20623
rect 410 20558 453 20622
rect 517 20558 560 20622
rect 23246 20558 23289 20622
rect 23353 20558 23396 20622
rect 452 20557 518 20558
rect 23288 20557 23354 20558
rect 452 20385 518 20386
rect 23288 20385 23354 20386
rect 410 20321 453 20385
rect 517 20321 560 20385
rect 23246 20321 23289 20385
rect 23353 20321 23396 20385
rect 452 20320 518 20321
rect 23288 20320 23354 20321
rect 452 20069 518 20070
rect 23288 20069 23354 20070
rect 410 20005 453 20069
rect 517 20005 560 20069
rect 23246 20005 23289 20069
rect 23353 20005 23396 20069
rect 452 20004 518 20005
rect 23288 20004 23354 20005
rect 452 19832 518 19833
rect 23288 19832 23354 19833
rect 410 19768 453 19832
rect 517 19768 560 19832
rect 23246 19768 23289 19832
rect 23353 19768 23396 19832
rect 452 19767 518 19768
rect 23288 19767 23354 19768
rect 452 19595 518 19596
rect 23288 19595 23354 19596
rect 410 19531 453 19595
rect 517 19531 560 19595
rect 23246 19531 23289 19595
rect 23353 19531 23396 19595
rect 452 19530 518 19531
rect 23288 19530 23354 19531
rect 452 19279 518 19280
rect 23288 19279 23354 19280
rect 410 19215 453 19279
rect 517 19215 560 19279
rect 23246 19215 23289 19279
rect 23353 19215 23396 19279
rect 452 19214 518 19215
rect 23288 19214 23354 19215
rect 452 19042 518 19043
rect 23288 19042 23354 19043
rect 410 18978 453 19042
rect 517 18978 560 19042
rect 23246 18978 23289 19042
rect 23353 18978 23396 19042
rect 452 18977 518 18978
rect 23288 18977 23354 18978
rect 452 18805 518 18806
rect 23288 18805 23354 18806
rect 410 18741 453 18805
rect 517 18741 560 18805
rect 23246 18741 23289 18805
rect 23353 18741 23396 18805
rect 452 18740 518 18741
rect 23288 18740 23354 18741
rect 452 18489 518 18490
rect 23288 18489 23354 18490
rect 410 18425 453 18489
rect 517 18425 560 18489
rect 23246 18425 23289 18489
rect 23353 18425 23396 18489
rect 452 18424 518 18425
rect 23288 18424 23354 18425
rect 452 18252 518 18253
rect 23288 18252 23354 18253
rect 410 18188 453 18252
rect 517 18188 560 18252
rect 23246 18188 23289 18252
rect 23353 18188 23396 18252
rect 452 18187 518 18188
rect 23288 18187 23354 18188
rect 452 18015 518 18016
rect 23288 18015 23354 18016
rect 410 17951 453 18015
rect 517 17951 560 18015
rect 23246 17951 23289 18015
rect 23353 17951 23396 18015
rect 452 17950 518 17951
rect 23288 17950 23354 17951
rect 452 17699 518 17700
rect 23288 17699 23354 17700
rect 410 17635 453 17699
rect 517 17635 560 17699
rect 23246 17635 23289 17699
rect 23353 17635 23396 17699
rect 452 17634 518 17635
rect 23288 17634 23354 17635
rect 452 17462 518 17463
rect 23288 17462 23354 17463
rect 410 17398 453 17462
rect 517 17398 560 17462
rect 23246 17398 23289 17462
rect 23353 17398 23396 17462
rect 452 17397 518 17398
rect 23288 17397 23354 17398
rect 452 17225 518 17226
rect 23288 17225 23354 17226
rect 410 17161 453 17225
rect 517 17161 560 17225
rect 23246 17161 23289 17225
rect 23353 17161 23396 17225
rect 452 17160 518 17161
rect 23288 17160 23354 17161
rect 452 16909 518 16910
rect 23288 16909 23354 16910
rect 410 16845 453 16909
rect 517 16845 560 16909
rect 23246 16845 23289 16909
rect 23353 16845 23396 16909
rect 452 16844 518 16845
rect 23288 16844 23354 16845
rect 452 16672 518 16673
rect 23288 16672 23354 16673
rect 410 16608 453 16672
rect 517 16608 560 16672
rect 23246 16608 23289 16672
rect 23353 16608 23396 16672
rect 452 16607 518 16608
rect 23288 16607 23354 16608
rect 452 16435 518 16436
rect 23288 16435 23354 16436
rect 410 16371 453 16435
rect 517 16371 560 16435
rect 23246 16371 23289 16435
rect 23353 16371 23396 16435
rect 452 16370 518 16371
rect 23288 16370 23354 16371
rect 452 16119 518 16120
rect 23288 16119 23354 16120
rect 410 16055 453 16119
rect 517 16055 560 16119
rect 23246 16055 23289 16119
rect 23353 16055 23396 16119
rect 452 16054 518 16055
rect 23288 16054 23354 16055
rect 452 15882 518 15883
rect 23288 15882 23354 15883
rect 410 15818 453 15882
rect 517 15818 560 15882
rect 23246 15818 23289 15882
rect 23353 15818 23396 15882
rect 452 15817 518 15818
rect 23288 15817 23354 15818
rect 452 15645 518 15646
rect 23288 15645 23354 15646
rect 410 15581 453 15645
rect 517 15581 560 15645
rect 23246 15581 23289 15645
rect 23353 15581 23396 15645
rect 452 15580 518 15581
rect 23288 15580 23354 15581
rect 452 15329 518 15330
rect 23288 15329 23354 15330
rect 410 15265 453 15329
rect 517 15265 560 15329
rect 23246 15265 23289 15329
rect 23353 15265 23396 15329
rect 452 15264 518 15265
rect 23288 15264 23354 15265
rect 452 15092 518 15093
rect 23288 15092 23354 15093
rect 410 15028 453 15092
rect 517 15028 560 15092
rect 23246 15028 23289 15092
rect 23353 15028 23396 15092
rect 452 15027 518 15028
rect 23288 15027 23354 15028
rect 452 14855 518 14856
rect 23288 14855 23354 14856
rect 410 14791 453 14855
rect 517 14791 560 14855
rect 23246 14791 23289 14855
rect 23353 14791 23396 14855
rect 452 14790 518 14791
rect 23288 14790 23354 14791
rect 452 14539 518 14540
rect 23288 14539 23354 14540
rect 410 14475 453 14539
rect 517 14475 560 14539
rect 23246 14475 23289 14539
rect 23353 14475 23396 14539
rect 452 14474 518 14475
rect 23288 14474 23354 14475
rect 452 14302 518 14303
rect 23288 14302 23354 14303
rect 410 14238 453 14302
rect 517 14238 560 14302
rect 23246 14238 23289 14302
rect 23353 14238 23396 14302
rect 452 14237 518 14238
rect 23288 14237 23354 14238
rect 452 14065 518 14066
rect 23288 14065 23354 14066
rect 410 14001 453 14065
rect 517 14001 560 14065
rect 23246 14001 23289 14065
rect 23353 14001 23396 14065
rect 452 14000 518 14001
rect 23288 14000 23354 14001
rect 452 13749 518 13750
rect 23288 13749 23354 13750
rect 410 13685 453 13749
rect 517 13685 560 13749
rect 23246 13685 23289 13749
rect 23353 13685 23396 13749
rect 452 13684 518 13685
rect 23288 13684 23354 13685
rect 452 13512 518 13513
rect 23288 13512 23354 13513
rect 410 13448 453 13512
rect 517 13448 560 13512
rect 23246 13448 23289 13512
rect 23353 13448 23396 13512
rect 452 13447 518 13448
rect 23288 13447 23354 13448
rect 452 13275 518 13276
rect 23288 13275 23354 13276
rect 410 13211 453 13275
rect 517 13211 560 13275
rect 23246 13211 23289 13275
rect 23353 13211 23396 13275
rect 452 13210 518 13211
rect 23288 13210 23354 13211
rect 452 12959 518 12960
rect 23288 12959 23354 12960
rect 410 12895 453 12959
rect 517 12895 560 12959
rect 23246 12895 23289 12959
rect 23353 12895 23396 12959
rect 452 12894 518 12895
rect 23288 12894 23354 12895
rect 452 12722 518 12723
rect 23288 12722 23354 12723
rect 410 12658 453 12722
rect 517 12658 560 12722
rect 23246 12658 23289 12722
rect 23353 12658 23396 12722
rect 452 12657 518 12658
rect 23288 12657 23354 12658
rect 452 12485 518 12486
rect 23288 12485 23354 12486
rect 410 12421 453 12485
rect 517 12421 560 12485
rect 23246 12421 23289 12485
rect 23353 12421 23396 12485
rect 452 12420 518 12421
rect 23288 12420 23354 12421
rect 452 12169 518 12170
rect 23288 12169 23354 12170
rect 410 12105 453 12169
rect 517 12105 560 12169
rect 23246 12105 23289 12169
rect 23353 12105 23396 12169
rect 452 12104 518 12105
rect 23288 12104 23354 12105
rect 452 11932 518 11933
rect 23288 11932 23354 11933
rect 410 11868 453 11932
rect 517 11868 560 11932
rect 23246 11868 23289 11932
rect 23353 11868 23396 11932
rect 452 11867 518 11868
rect 23288 11867 23354 11868
rect 452 11695 518 11696
rect 23288 11695 23354 11696
rect 410 11631 453 11695
rect 517 11631 560 11695
rect 23246 11631 23289 11695
rect 23353 11631 23396 11695
rect 452 11630 518 11631
rect 23288 11630 23354 11631
rect 452 11379 518 11380
rect 23288 11379 23354 11380
rect 410 11315 453 11379
rect 517 11315 560 11379
rect 23246 11315 23289 11379
rect 23353 11315 23396 11379
rect 452 11314 518 11315
rect 23288 11314 23354 11315
rect 452 11142 518 11143
rect 23288 11142 23354 11143
rect 410 11078 453 11142
rect 517 11078 560 11142
rect 23246 11078 23289 11142
rect 23353 11078 23396 11142
rect 452 11077 518 11078
rect 23288 11077 23354 11078
rect 452 10905 518 10906
rect 23288 10905 23354 10906
rect 410 10841 453 10905
rect 517 10841 560 10905
rect 23246 10841 23289 10905
rect 23353 10841 23396 10905
rect 452 10840 518 10841
rect 23288 10840 23354 10841
rect 452 10589 518 10590
rect 23288 10589 23354 10590
rect 410 10525 453 10589
rect 517 10525 560 10589
rect 23246 10525 23289 10589
rect 23353 10525 23396 10589
rect 452 10524 518 10525
rect 23288 10524 23354 10525
rect 452 10352 518 10353
rect 23288 10352 23354 10353
rect 410 10288 453 10352
rect 517 10288 560 10352
rect 23246 10288 23289 10352
rect 23353 10288 23396 10352
rect 452 10287 518 10288
rect 23288 10287 23354 10288
rect 452 10115 518 10116
rect 23288 10115 23354 10116
rect 410 10051 453 10115
rect 517 10051 560 10115
rect 23246 10051 23289 10115
rect 23353 10051 23396 10115
rect 452 10050 518 10051
rect 23288 10050 23354 10051
rect 452 9799 518 9800
rect 23288 9799 23354 9800
rect 410 9735 453 9799
rect 517 9735 560 9799
rect 23246 9735 23289 9799
rect 23353 9735 23396 9799
rect 452 9734 518 9735
rect 23288 9734 23354 9735
rect 452 9562 518 9563
rect 23288 9562 23354 9563
rect 410 9498 453 9562
rect 517 9498 560 9562
rect 23246 9498 23289 9562
rect 23353 9498 23396 9562
rect 452 9497 518 9498
rect 23288 9497 23354 9498
rect 452 9325 518 9326
rect 23288 9325 23354 9326
rect 410 9261 453 9325
rect 517 9261 560 9325
rect 23246 9261 23289 9325
rect 23353 9261 23396 9325
rect 452 9260 518 9261
rect 23288 9260 23354 9261
rect 452 9009 518 9010
rect 23288 9009 23354 9010
rect 410 8945 453 9009
rect 517 8945 560 9009
rect 23246 8945 23289 9009
rect 23353 8945 23396 9009
rect 452 8944 518 8945
rect 23288 8944 23354 8945
rect 452 8772 518 8773
rect 23288 8772 23354 8773
rect 410 8708 453 8772
rect 517 8708 560 8772
rect 23246 8708 23289 8772
rect 23353 8708 23396 8772
rect 452 8707 518 8708
rect 23288 8707 23354 8708
rect 452 8535 518 8536
rect 23288 8535 23354 8536
rect 410 8471 453 8535
rect 517 8471 560 8535
rect 23246 8471 23289 8535
rect 23353 8471 23396 8535
rect 452 8470 518 8471
rect 23288 8470 23354 8471
rect 452 8219 518 8220
rect 23288 8219 23354 8220
rect 410 8155 453 8219
rect 517 8155 560 8219
rect 23246 8155 23289 8219
rect 23353 8155 23396 8219
rect 452 8154 518 8155
rect 23288 8154 23354 8155
rect 452 7982 518 7983
rect 23288 7982 23354 7983
rect 410 7918 453 7982
rect 517 7918 560 7982
rect 23246 7918 23289 7982
rect 23353 7918 23396 7982
rect 452 7917 518 7918
rect 23288 7917 23354 7918
rect 452 7745 518 7746
rect 23288 7745 23354 7746
rect 410 7681 453 7745
rect 517 7681 560 7745
rect 23246 7681 23289 7745
rect 23353 7681 23396 7745
rect 452 7680 518 7681
rect 23288 7680 23354 7681
rect 452 7429 518 7430
rect 23288 7429 23354 7430
rect 410 7365 453 7429
rect 517 7365 560 7429
rect 23246 7365 23289 7429
rect 23353 7365 23396 7429
rect 452 7364 518 7365
rect 23288 7364 23354 7365
rect 452 7192 518 7193
rect 23288 7192 23354 7193
rect 410 7128 453 7192
rect 517 7128 560 7192
rect 23246 7128 23289 7192
rect 23353 7128 23396 7192
rect 452 7127 518 7128
rect 23288 7127 23354 7128
rect 452 6955 518 6956
rect 23288 6955 23354 6956
rect 410 6891 453 6955
rect 517 6891 560 6955
rect 23246 6891 23289 6955
rect 23353 6891 23396 6955
rect 452 6890 518 6891
rect 23288 6890 23354 6891
rect 452 6639 518 6640
rect 23288 6639 23354 6640
rect 410 6575 453 6639
rect 517 6575 560 6639
rect 23246 6575 23289 6639
rect 23353 6575 23396 6639
rect 452 6574 518 6575
rect 23288 6574 23354 6575
rect 452 6402 518 6403
rect 23288 6402 23354 6403
rect 410 6338 453 6402
rect 517 6338 560 6402
rect 23246 6338 23289 6402
rect 23353 6338 23396 6402
rect 452 6337 518 6338
rect 23288 6337 23354 6338
rect 452 6165 518 6166
rect 23288 6165 23354 6166
rect 410 6101 453 6165
rect 517 6101 560 6165
rect 23246 6101 23289 6165
rect 23353 6101 23396 6165
rect 452 6100 518 6101
rect 23288 6100 23354 6101
rect 452 5849 518 5850
rect 23288 5849 23354 5850
rect 410 5785 453 5849
rect 517 5785 560 5849
rect 23246 5785 23289 5849
rect 23353 5785 23396 5849
rect 452 5784 518 5785
rect 23288 5784 23354 5785
rect 452 5612 518 5613
rect 23288 5612 23354 5613
rect 410 5548 453 5612
rect 517 5548 560 5612
rect 23246 5548 23289 5612
rect 23353 5548 23396 5612
rect 452 5547 518 5548
rect 23288 5547 23354 5548
rect 452 5375 518 5376
rect 23288 5375 23354 5376
rect 410 5311 453 5375
rect 517 5311 560 5375
rect 23246 5311 23289 5375
rect 23353 5311 23396 5375
rect 452 5310 518 5311
rect 23288 5310 23354 5311
rect 452 5059 518 5060
rect 23288 5059 23354 5060
rect 410 4995 453 5059
rect 517 4995 560 5059
rect 23246 4995 23289 5059
rect 23353 4995 23396 5059
rect 452 4994 518 4995
rect 23288 4994 23354 4995
rect 452 4822 518 4823
rect 23288 4822 23354 4823
rect 410 4758 453 4822
rect 517 4758 560 4822
rect 23246 4758 23289 4822
rect 23353 4758 23396 4822
rect 452 4757 518 4758
rect 23288 4757 23354 4758
rect 452 4585 518 4586
rect 23288 4585 23354 4586
rect 410 4521 453 4585
rect 517 4521 560 4585
rect 23246 4521 23289 4585
rect 23353 4521 23396 4585
rect 452 4520 518 4521
rect 23288 4520 23354 4521
rect 452 4269 518 4270
rect 23288 4269 23354 4270
rect 410 4205 453 4269
rect 517 4205 560 4269
rect 23246 4205 23289 4269
rect 23353 4205 23396 4269
rect 452 4204 518 4205
rect 23288 4204 23354 4205
rect 452 4032 518 4033
rect 23288 4032 23354 4033
rect 410 3968 453 4032
rect 517 3968 560 4032
rect 23246 3968 23289 4032
rect 23353 3968 23396 4032
rect 452 3967 518 3968
rect 23288 3967 23354 3968
rect 452 3795 518 3796
rect 23288 3795 23354 3796
rect 410 3731 453 3795
rect 517 3731 560 3795
rect 23246 3731 23289 3795
rect 23353 3731 23396 3795
rect 452 3730 518 3731
rect 23288 3730 23354 3731
rect 452 3479 518 3480
rect 23288 3479 23354 3480
rect 410 3415 453 3479
rect 517 3415 560 3479
rect 23246 3415 23289 3479
rect 23353 3415 23396 3479
rect 452 3414 518 3415
rect 23288 3414 23354 3415
rect 452 3242 518 3243
rect 23288 3242 23354 3243
rect 410 3178 453 3242
rect 517 3178 560 3242
rect 23246 3178 23289 3242
rect 23353 3178 23396 3242
rect 452 3177 518 3178
rect 23288 3177 23354 3178
rect 452 3005 518 3006
rect 23288 3005 23354 3006
rect 410 2941 453 3005
rect 517 2941 560 3005
rect 23246 2941 23289 3005
rect 23353 2941 23396 3005
rect 452 2940 518 2941
rect 23288 2940 23354 2941
rect 452 2689 518 2690
rect 23288 2689 23354 2690
rect 410 2625 453 2689
rect 517 2625 560 2689
rect 23246 2625 23289 2689
rect 23353 2625 23396 2689
rect 452 2624 518 2625
rect 23288 2624 23354 2625
rect 452 2452 518 2453
rect 23288 2452 23354 2453
rect 410 2388 453 2452
rect 517 2388 560 2452
rect 23246 2388 23289 2452
rect 23353 2388 23396 2452
rect 452 2387 518 2388
rect 23288 2387 23354 2388
rect 452 2215 518 2216
rect 23288 2215 23354 2216
rect 410 2151 453 2215
rect 517 2151 560 2215
rect 23246 2151 23289 2215
rect 23353 2151 23396 2215
rect 452 2150 518 2151
rect 23288 2150 23354 2151
rect 452 1899 518 1900
rect 23288 1899 23354 1900
rect 410 1835 453 1899
rect 517 1835 560 1899
rect 23246 1835 23289 1899
rect 23353 1835 23396 1899
rect 452 1834 518 1835
rect 23288 1834 23354 1835
rect 452 1662 518 1663
rect 23288 1662 23354 1663
rect 410 1598 453 1662
rect 517 1598 560 1662
rect 23246 1598 23289 1662
rect 23353 1598 23396 1662
rect 452 1597 518 1598
rect 23288 1597 23354 1598
rect 452 1425 518 1426
rect 23288 1425 23354 1426
rect 410 1361 453 1425
rect 517 1361 560 1425
rect 23246 1361 23289 1425
rect 23353 1361 23396 1425
rect 452 1360 518 1361
rect 23288 1360 23354 1361
rect 452 1109 518 1110
rect 23288 1109 23354 1110
rect 410 1045 453 1109
rect 517 1045 560 1109
rect 23246 1045 23289 1109
rect 23353 1045 23396 1109
rect 452 1044 518 1045
rect 23288 1044 23354 1045
rect 452 872 518 873
rect 23288 872 23354 873
rect 410 808 453 872
rect 517 808 560 872
rect 23246 808 23289 872
rect 23353 808 23396 872
rect 452 807 518 808
rect 23288 807 23354 808
rect 452 745 518 746
rect 23288 745 23354 746
rect 410 681 453 745
rect 517 681 560 745
rect 23246 681 23289 745
rect 23353 681 23396 745
rect 452 680 518 681
rect 23288 680 23354 681
rect 42 311 108 312
rect 23698 311 23764 312
rect 0 247 43 311
rect 107 247 150 311
rect 23656 247 23699 311
rect 23763 247 23806 311
rect 42 246 108 247
rect 23698 246 23764 247
<< via3 >>
rect 43 26709 107 26713
rect 43 26653 47 26709
rect 47 26653 103 26709
rect 103 26653 107 26709
rect 43 26649 107 26653
rect 23699 26709 23763 26713
rect 23699 26653 23703 26709
rect 23703 26653 23759 26709
rect 23759 26653 23763 26709
rect 23699 26649 23763 26653
rect 453 26495 517 26499
rect 453 26439 457 26495
rect 457 26439 513 26495
rect 513 26439 517 26495
rect 453 26435 517 26439
rect 23289 26495 23353 26499
rect 23289 26439 23293 26495
rect 23293 26439 23349 26495
rect 23349 26439 23353 26495
rect 23289 26435 23353 26439
rect 453 26148 517 26152
rect 453 26092 457 26148
rect 457 26092 513 26148
rect 513 26092 517 26148
rect 453 26088 517 26092
rect 23289 26148 23353 26152
rect 23289 26092 23293 26148
rect 23293 26092 23349 26148
rect 23349 26092 23353 26148
rect 23289 26088 23353 26092
rect 453 25911 517 25915
rect 453 25855 457 25911
rect 457 25855 513 25911
rect 513 25855 517 25911
rect 453 25851 517 25855
rect 23289 25911 23353 25915
rect 23289 25855 23293 25911
rect 23293 25855 23349 25911
rect 23349 25855 23353 25911
rect 23289 25851 23353 25855
rect 453 25595 517 25599
rect 453 25539 457 25595
rect 457 25539 513 25595
rect 513 25539 517 25595
rect 453 25535 517 25539
rect 23289 25595 23353 25599
rect 23289 25539 23293 25595
rect 23293 25539 23349 25595
rect 23349 25539 23353 25595
rect 23289 25535 23353 25539
rect 453 25358 517 25362
rect 453 25302 457 25358
rect 457 25302 513 25358
rect 513 25302 517 25358
rect 453 25298 517 25302
rect 23289 25358 23353 25362
rect 23289 25302 23293 25358
rect 23293 25302 23349 25358
rect 23349 25302 23353 25358
rect 23289 25298 23353 25302
rect 453 25121 517 25125
rect 453 25065 457 25121
rect 457 25065 513 25121
rect 513 25065 517 25121
rect 453 25061 517 25065
rect 23289 25121 23353 25125
rect 23289 25065 23293 25121
rect 23293 25065 23349 25121
rect 23349 25065 23353 25121
rect 23289 25061 23353 25065
rect 453 24805 517 24809
rect 453 24749 457 24805
rect 457 24749 513 24805
rect 513 24749 517 24805
rect 453 24745 517 24749
rect 23289 24805 23353 24809
rect 23289 24749 23293 24805
rect 23293 24749 23349 24805
rect 23349 24749 23353 24805
rect 23289 24745 23353 24749
rect 453 24568 517 24572
rect 453 24512 457 24568
rect 457 24512 513 24568
rect 513 24512 517 24568
rect 453 24508 517 24512
rect 23289 24568 23353 24572
rect 23289 24512 23293 24568
rect 23293 24512 23349 24568
rect 23349 24512 23353 24568
rect 23289 24508 23353 24512
rect 453 24331 517 24335
rect 453 24275 457 24331
rect 457 24275 513 24331
rect 513 24275 517 24331
rect 453 24271 517 24275
rect 23289 24331 23353 24335
rect 23289 24275 23293 24331
rect 23293 24275 23349 24331
rect 23349 24275 23353 24331
rect 23289 24271 23353 24275
rect 453 24015 517 24019
rect 453 23959 457 24015
rect 457 23959 513 24015
rect 513 23959 517 24015
rect 453 23955 517 23959
rect 23289 24015 23353 24019
rect 23289 23959 23293 24015
rect 23293 23959 23349 24015
rect 23349 23959 23353 24015
rect 23289 23955 23353 23959
rect 453 23778 517 23782
rect 453 23722 457 23778
rect 457 23722 513 23778
rect 513 23722 517 23778
rect 453 23718 517 23722
rect 23289 23778 23353 23782
rect 23289 23722 23293 23778
rect 23293 23722 23349 23778
rect 23349 23722 23353 23778
rect 23289 23718 23353 23722
rect 453 23541 517 23545
rect 453 23485 457 23541
rect 457 23485 513 23541
rect 513 23485 517 23541
rect 453 23481 517 23485
rect 23289 23541 23353 23545
rect 23289 23485 23293 23541
rect 23293 23485 23349 23541
rect 23349 23485 23353 23541
rect 23289 23481 23353 23485
rect 453 23225 517 23229
rect 453 23169 457 23225
rect 457 23169 513 23225
rect 513 23169 517 23225
rect 453 23165 517 23169
rect 23289 23225 23353 23229
rect 23289 23169 23293 23225
rect 23293 23169 23349 23225
rect 23349 23169 23353 23225
rect 23289 23165 23353 23169
rect 453 22988 517 22992
rect 453 22932 457 22988
rect 457 22932 513 22988
rect 513 22932 517 22988
rect 453 22928 517 22932
rect 23289 22988 23353 22992
rect 23289 22932 23293 22988
rect 23293 22932 23349 22988
rect 23349 22932 23353 22988
rect 23289 22928 23353 22932
rect 453 22751 517 22755
rect 453 22695 457 22751
rect 457 22695 513 22751
rect 513 22695 517 22751
rect 453 22691 517 22695
rect 23289 22751 23353 22755
rect 23289 22695 23293 22751
rect 23293 22695 23349 22751
rect 23349 22695 23353 22751
rect 23289 22691 23353 22695
rect 453 22435 517 22439
rect 453 22379 457 22435
rect 457 22379 513 22435
rect 513 22379 517 22435
rect 453 22375 517 22379
rect 23289 22435 23353 22439
rect 23289 22379 23293 22435
rect 23293 22379 23349 22435
rect 23349 22379 23353 22435
rect 23289 22375 23353 22379
rect 453 22198 517 22202
rect 453 22142 457 22198
rect 457 22142 513 22198
rect 513 22142 517 22198
rect 453 22138 517 22142
rect 23289 22198 23353 22202
rect 23289 22142 23293 22198
rect 23293 22142 23349 22198
rect 23349 22142 23353 22198
rect 23289 22138 23353 22142
rect 453 21961 517 21965
rect 453 21905 457 21961
rect 457 21905 513 21961
rect 513 21905 517 21961
rect 453 21901 517 21905
rect 23289 21961 23353 21965
rect 23289 21905 23293 21961
rect 23293 21905 23349 21961
rect 23349 21905 23353 21961
rect 23289 21901 23353 21905
rect 453 21645 517 21649
rect 453 21589 457 21645
rect 457 21589 513 21645
rect 513 21589 517 21645
rect 453 21585 517 21589
rect 23289 21645 23353 21649
rect 23289 21589 23293 21645
rect 23293 21589 23349 21645
rect 23349 21589 23353 21645
rect 23289 21585 23353 21589
rect 453 21408 517 21412
rect 453 21352 457 21408
rect 457 21352 513 21408
rect 513 21352 517 21408
rect 453 21348 517 21352
rect 23289 21408 23353 21412
rect 23289 21352 23293 21408
rect 23293 21352 23349 21408
rect 23349 21352 23353 21408
rect 23289 21348 23353 21352
rect 453 21171 517 21175
rect 453 21115 457 21171
rect 457 21115 513 21171
rect 513 21115 517 21171
rect 453 21111 517 21115
rect 23289 21171 23353 21175
rect 23289 21115 23293 21171
rect 23293 21115 23349 21171
rect 23349 21115 23353 21171
rect 23289 21111 23353 21115
rect 453 20855 517 20859
rect 453 20799 457 20855
rect 457 20799 513 20855
rect 513 20799 517 20855
rect 453 20795 517 20799
rect 23289 20855 23353 20859
rect 23289 20799 23293 20855
rect 23293 20799 23349 20855
rect 23349 20799 23353 20855
rect 23289 20795 23353 20799
rect 453 20618 517 20622
rect 453 20562 457 20618
rect 457 20562 513 20618
rect 513 20562 517 20618
rect 453 20558 517 20562
rect 23289 20618 23353 20622
rect 23289 20562 23293 20618
rect 23293 20562 23349 20618
rect 23349 20562 23353 20618
rect 23289 20558 23353 20562
rect 453 20381 517 20385
rect 453 20325 457 20381
rect 457 20325 513 20381
rect 513 20325 517 20381
rect 453 20321 517 20325
rect 23289 20381 23353 20385
rect 23289 20325 23293 20381
rect 23293 20325 23349 20381
rect 23349 20325 23353 20381
rect 23289 20321 23353 20325
rect 453 20065 517 20069
rect 453 20009 457 20065
rect 457 20009 513 20065
rect 513 20009 517 20065
rect 453 20005 517 20009
rect 23289 20065 23353 20069
rect 23289 20009 23293 20065
rect 23293 20009 23349 20065
rect 23349 20009 23353 20065
rect 23289 20005 23353 20009
rect 453 19828 517 19832
rect 453 19772 457 19828
rect 457 19772 513 19828
rect 513 19772 517 19828
rect 453 19768 517 19772
rect 23289 19828 23353 19832
rect 23289 19772 23293 19828
rect 23293 19772 23349 19828
rect 23349 19772 23353 19828
rect 23289 19768 23353 19772
rect 453 19591 517 19595
rect 453 19535 457 19591
rect 457 19535 513 19591
rect 513 19535 517 19591
rect 453 19531 517 19535
rect 23289 19591 23353 19595
rect 23289 19535 23293 19591
rect 23293 19535 23349 19591
rect 23349 19535 23353 19591
rect 23289 19531 23353 19535
rect 453 19275 517 19279
rect 453 19219 457 19275
rect 457 19219 513 19275
rect 513 19219 517 19275
rect 453 19215 517 19219
rect 23289 19275 23353 19279
rect 23289 19219 23293 19275
rect 23293 19219 23349 19275
rect 23349 19219 23353 19275
rect 23289 19215 23353 19219
rect 453 19038 517 19042
rect 453 18982 457 19038
rect 457 18982 513 19038
rect 513 18982 517 19038
rect 453 18978 517 18982
rect 23289 19038 23353 19042
rect 23289 18982 23293 19038
rect 23293 18982 23349 19038
rect 23349 18982 23353 19038
rect 23289 18978 23353 18982
rect 453 18801 517 18805
rect 453 18745 457 18801
rect 457 18745 513 18801
rect 513 18745 517 18801
rect 453 18741 517 18745
rect 23289 18801 23353 18805
rect 23289 18745 23293 18801
rect 23293 18745 23349 18801
rect 23349 18745 23353 18801
rect 23289 18741 23353 18745
rect 453 18485 517 18489
rect 453 18429 457 18485
rect 457 18429 513 18485
rect 513 18429 517 18485
rect 453 18425 517 18429
rect 23289 18485 23353 18489
rect 23289 18429 23293 18485
rect 23293 18429 23349 18485
rect 23349 18429 23353 18485
rect 23289 18425 23353 18429
rect 453 18248 517 18252
rect 453 18192 457 18248
rect 457 18192 513 18248
rect 513 18192 517 18248
rect 453 18188 517 18192
rect 23289 18248 23353 18252
rect 23289 18192 23293 18248
rect 23293 18192 23349 18248
rect 23349 18192 23353 18248
rect 23289 18188 23353 18192
rect 453 18011 517 18015
rect 453 17955 457 18011
rect 457 17955 513 18011
rect 513 17955 517 18011
rect 453 17951 517 17955
rect 23289 18011 23353 18015
rect 23289 17955 23293 18011
rect 23293 17955 23349 18011
rect 23349 17955 23353 18011
rect 23289 17951 23353 17955
rect 453 17695 517 17699
rect 453 17639 457 17695
rect 457 17639 513 17695
rect 513 17639 517 17695
rect 453 17635 517 17639
rect 23289 17695 23353 17699
rect 23289 17639 23293 17695
rect 23293 17639 23349 17695
rect 23349 17639 23353 17695
rect 23289 17635 23353 17639
rect 453 17458 517 17462
rect 453 17402 457 17458
rect 457 17402 513 17458
rect 513 17402 517 17458
rect 453 17398 517 17402
rect 23289 17458 23353 17462
rect 23289 17402 23293 17458
rect 23293 17402 23349 17458
rect 23349 17402 23353 17458
rect 23289 17398 23353 17402
rect 453 17221 517 17225
rect 453 17165 457 17221
rect 457 17165 513 17221
rect 513 17165 517 17221
rect 453 17161 517 17165
rect 23289 17221 23353 17225
rect 23289 17165 23293 17221
rect 23293 17165 23349 17221
rect 23349 17165 23353 17221
rect 23289 17161 23353 17165
rect 453 16905 517 16909
rect 453 16849 457 16905
rect 457 16849 513 16905
rect 513 16849 517 16905
rect 453 16845 517 16849
rect 23289 16905 23353 16909
rect 23289 16849 23293 16905
rect 23293 16849 23349 16905
rect 23349 16849 23353 16905
rect 23289 16845 23353 16849
rect 453 16668 517 16672
rect 453 16612 457 16668
rect 457 16612 513 16668
rect 513 16612 517 16668
rect 453 16608 517 16612
rect 23289 16668 23353 16672
rect 23289 16612 23293 16668
rect 23293 16612 23349 16668
rect 23349 16612 23353 16668
rect 23289 16608 23353 16612
rect 453 16431 517 16435
rect 453 16375 457 16431
rect 457 16375 513 16431
rect 513 16375 517 16431
rect 453 16371 517 16375
rect 23289 16431 23353 16435
rect 23289 16375 23293 16431
rect 23293 16375 23349 16431
rect 23349 16375 23353 16431
rect 23289 16371 23353 16375
rect 453 16115 517 16119
rect 453 16059 457 16115
rect 457 16059 513 16115
rect 513 16059 517 16115
rect 453 16055 517 16059
rect 23289 16115 23353 16119
rect 23289 16059 23293 16115
rect 23293 16059 23349 16115
rect 23349 16059 23353 16115
rect 23289 16055 23353 16059
rect 453 15878 517 15882
rect 453 15822 457 15878
rect 457 15822 513 15878
rect 513 15822 517 15878
rect 453 15818 517 15822
rect 23289 15878 23353 15882
rect 23289 15822 23293 15878
rect 23293 15822 23349 15878
rect 23349 15822 23353 15878
rect 23289 15818 23353 15822
rect 453 15641 517 15645
rect 453 15585 457 15641
rect 457 15585 513 15641
rect 513 15585 517 15641
rect 453 15581 517 15585
rect 23289 15641 23353 15645
rect 23289 15585 23293 15641
rect 23293 15585 23349 15641
rect 23349 15585 23353 15641
rect 23289 15581 23353 15585
rect 453 15325 517 15329
rect 453 15269 457 15325
rect 457 15269 513 15325
rect 513 15269 517 15325
rect 453 15265 517 15269
rect 23289 15325 23353 15329
rect 23289 15269 23293 15325
rect 23293 15269 23349 15325
rect 23349 15269 23353 15325
rect 23289 15265 23353 15269
rect 453 15088 517 15092
rect 453 15032 457 15088
rect 457 15032 513 15088
rect 513 15032 517 15088
rect 453 15028 517 15032
rect 23289 15088 23353 15092
rect 23289 15032 23293 15088
rect 23293 15032 23349 15088
rect 23349 15032 23353 15088
rect 23289 15028 23353 15032
rect 453 14851 517 14855
rect 453 14795 457 14851
rect 457 14795 513 14851
rect 513 14795 517 14851
rect 453 14791 517 14795
rect 23289 14851 23353 14855
rect 23289 14795 23293 14851
rect 23293 14795 23349 14851
rect 23349 14795 23353 14851
rect 23289 14791 23353 14795
rect 453 14535 517 14539
rect 453 14479 457 14535
rect 457 14479 513 14535
rect 513 14479 517 14535
rect 453 14475 517 14479
rect 23289 14535 23353 14539
rect 23289 14479 23293 14535
rect 23293 14479 23349 14535
rect 23349 14479 23353 14535
rect 23289 14475 23353 14479
rect 453 14298 517 14302
rect 453 14242 457 14298
rect 457 14242 513 14298
rect 513 14242 517 14298
rect 453 14238 517 14242
rect 23289 14298 23353 14302
rect 23289 14242 23293 14298
rect 23293 14242 23349 14298
rect 23349 14242 23353 14298
rect 23289 14238 23353 14242
rect 453 14061 517 14065
rect 453 14005 457 14061
rect 457 14005 513 14061
rect 513 14005 517 14061
rect 453 14001 517 14005
rect 23289 14061 23353 14065
rect 23289 14005 23293 14061
rect 23293 14005 23349 14061
rect 23349 14005 23353 14061
rect 23289 14001 23353 14005
rect 453 13745 517 13749
rect 453 13689 457 13745
rect 457 13689 513 13745
rect 513 13689 517 13745
rect 453 13685 517 13689
rect 23289 13745 23353 13749
rect 23289 13689 23293 13745
rect 23293 13689 23349 13745
rect 23349 13689 23353 13745
rect 23289 13685 23353 13689
rect 453 13508 517 13512
rect 453 13452 457 13508
rect 457 13452 513 13508
rect 513 13452 517 13508
rect 453 13448 517 13452
rect 23289 13508 23353 13512
rect 23289 13452 23293 13508
rect 23293 13452 23349 13508
rect 23349 13452 23353 13508
rect 23289 13448 23353 13452
rect 453 13271 517 13275
rect 453 13215 457 13271
rect 457 13215 513 13271
rect 513 13215 517 13271
rect 453 13211 517 13215
rect 23289 13271 23353 13275
rect 23289 13215 23293 13271
rect 23293 13215 23349 13271
rect 23349 13215 23353 13271
rect 23289 13211 23353 13215
rect 453 12955 517 12959
rect 453 12899 457 12955
rect 457 12899 513 12955
rect 513 12899 517 12955
rect 453 12895 517 12899
rect 23289 12955 23353 12959
rect 23289 12899 23293 12955
rect 23293 12899 23349 12955
rect 23349 12899 23353 12955
rect 23289 12895 23353 12899
rect 453 12718 517 12722
rect 453 12662 457 12718
rect 457 12662 513 12718
rect 513 12662 517 12718
rect 453 12658 517 12662
rect 23289 12718 23353 12722
rect 23289 12662 23293 12718
rect 23293 12662 23349 12718
rect 23349 12662 23353 12718
rect 23289 12658 23353 12662
rect 453 12481 517 12485
rect 453 12425 457 12481
rect 457 12425 513 12481
rect 513 12425 517 12481
rect 453 12421 517 12425
rect 23289 12481 23353 12485
rect 23289 12425 23293 12481
rect 23293 12425 23349 12481
rect 23349 12425 23353 12481
rect 23289 12421 23353 12425
rect 453 12165 517 12169
rect 453 12109 457 12165
rect 457 12109 513 12165
rect 513 12109 517 12165
rect 453 12105 517 12109
rect 23289 12165 23353 12169
rect 23289 12109 23293 12165
rect 23293 12109 23349 12165
rect 23349 12109 23353 12165
rect 23289 12105 23353 12109
rect 453 11928 517 11932
rect 453 11872 457 11928
rect 457 11872 513 11928
rect 513 11872 517 11928
rect 453 11868 517 11872
rect 23289 11928 23353 11932
rect 23289 11872 23293 11928
rect 23293 11872 23349 11928
rect 23349 11872 23353 11928
rect 23289 11868 23353 11872
rect 453 11691 517 11695
rect 453 11635 457 11691
rect 457 11635 513 11691
rect 513 11635 517 11691
rect 453 11631 517 11635
rect 23289 11691 23353 11695
rect 23289 11635 23293 11691
rect 23293 11635 23349 11691
rect 23349 11635 23353 11691
rect 23289 11631 23353 11635
rect 453 11375 517 11379
rect 453 11319 457 11375
rect 457 11319 513 11375
rect 513 11319 517 11375
rect 453 11315 517 11319
rect 23289 11375 23353 11379
rect 23289 11319 23293 11375
rect 23293 11319 23349 11375
rect 23349 11319 23353 11375
rect 23289 11315 23353 11319
rect 453 11138 517 11142
rect 453 11082 457 11138
rect 457 11082 513 11138
rect 513 11082 517 11138
rect 453 11078 517 11082
rect 23289 11138 23353 11142
rect 23289 11082 23293 11138
rect 23293 11082 23349 11138
rect 23349 11082 23353 11138
rect 23289 11078 23353 11082
rect 453 10901 517 10905
rect 453 10845 457 10901
rect 457 10845 513 10901
rect 513 10845 517 10901
rect 453 10841 517 10845
rect 23289 10901 23353 10905
rect 23289 10845 23293 10901
rect 23293 10845 23349 10901
rect 23349 10845 23353 10901
rect 23289 10841 23353 10845
rect 453 10585 517 10589
rect 453 10529 457 10585
rect 457 10529 513 10585
rect 513 10529 517 10585
rect 453 10525 517 10529
rect 23289 10585 23353 10589
rect 23289 10529 23293 10585
rect 23293 10529 23349 10585
rect 23349 10529 23353 10585
rect 23289 10525 23353 10529
rect 453 10348 517 10352
rect 453 10292 457 10348
rect 457 10292 513 10348
rect 513 10292 517 10348
rect 453 10288 517 10292
rect 23289 10348 23353 10352
rect 23289 10292 23293 10348
rect 23293 10292 23349 10348
rect 23349 10292 23353 10348
rect 23289 10288 23353 10292
rect 453 10111 517 10115
rect 453 10055 457 10111
rect 457 10055 513 10111
rect 513 10055 517 10111
rect 453 10051 517 10055
rect 23289 10111 23353 10115
rect 23289 10055 23293 10111
rect 23293 10055 23349 10111
rect 23349 10055 23353 10111
rect 23289 10051 23353 10055
rect 453 9795 517 9799
rect 453 9739 457 9795
rect 457 9739 513 9795
rect 513 9739 517 9795
rect 453 9735 517 9739
rect 23289 9795 23353 9799
rect 23289 9739 23293 9795
rect 23293 9739 23349 9795
rect 23349 9739 23353 9795
rect 23289 9735 23353 9739
rect 453 9558 517 9562
rect 453 9502 457 9558
rect 457 9502 513 9558
rect 513 9502 517 9558
rect 453 9498 517 9502
rect 23289 9558 23353 9562
rect 23289 9502 23293 9558
rect 23293 9502 23349 9558
rect 23349 9502 23353 9558
rect 23289 9498 23353 9502
rect 453 9321 517 9325
rect 453 9265 457 9321
rect 457 9265 513 9321
rect 513 9265 517 9321
rect 453 9261 517 9265
rect 23289 9321 23353 9325
rect 23289 9265 23293 9321
rect 23293 9265 23349 9321
rect 23349 9265 23353 9321
rect 23289 9261 23353 9265
rect 453 9005 517 9009
rect 453 8949 457 9005
rect 457 8949 513 9005
rect 513 8949 517 9005
rect 453 8945 517 8949
rect 23289 9005 23353 9009
rect 23289 8949 23293 9005
rect 23293 8949 23349 9005
rect 23349 8949 23353 9005
rect 23289 8945 23353 8949
rect 453 8768 517 8772
rect 453 8712 457 8768
rect 457 8712 513 8768
rect 513 8712 517 8768
rect 453 8708 517 8712
rect 23289 8768 23353 8772
rect 23289 8712 23293 8768
rect 23293 8712 23349 8768
rect 23349 8712 23353 8768
rect 23289 8708 23353 8712
rect 453 8531 517 8535
rect 453 8475 457 8531
rect 457 8475 513 8531
rect 513 8475 517 8531
rect 453 8471 517 8475
rect 23289 8531 23353 8535
rect 23289 8475 23293 8531
rect 23293 8475 23349 8531
rect 23349 8475 23353 8531
rect 23289 8471 23353 8475
rect 453 8215 517 8219
rect 453 8159 457 8215
rect 457 8159 513 8215
rect 513 8159 517 8215
rect 453 8155 517 8159
rect 23289 8215 23353 8219
rect 23289 8159 23293 8215
rect 23293 8159 23349 8215
rect 23349 8159 23353 8215
rect 23289 8155 23353 8159
rect 453 7978 517 7982
rect 453 7922 457 7978
rect 457 7922 513 7978
rect 513 7922 517 7978
rect 453 7918 517 7922
rect 23289 7978 23353 7982
rect 23289 7922 23293 7978
rect 23293 7922 23349 7978
rect 23349 7922 23353 7978
rect 23289 7918 23353 7922
rect 453 7741 517 7745
rect 453 7685 457 7741
rect 457 7685 513 7741
rect 513 7685 517 7741
rect 453 7681 517 7685
rect 23289 7741 23353 7745
rect 23289 7685 23293 7741
rect 23293 7685 23349 7741
rect 23349 7685 23353 7741
rect 23289 7681 23353 7685
rect 453 7425 517 7429
rect 453 7369 457 7425
rect 457 7369 513 7425
rect 513 7369 517 7425
rect 453 7365 517 7369
rect 23289 7425 23353 7429
rect 23289 7369 23293 7425
rect 23293 7369 23349 7425
rect 23349 7369 23353 7425
rect 23289 7365 23353 7369
rect 453 7188 517 7192
rect 453 7132 457 7188
rect 457 7132 513 7188
rect 513 7132 517 7188
rect 453 7128 517 7132
rect 23289 7188 23353 7192
rect 23289 7132 23293 7188
rect 23293 7132 23349 7188
rect 23349 7132 23353 7188
rect 23289 7128 23353 7132
rect 453 6951 517 6955
rect 453 6895 457 6951
rect 457 6895 513 6951
rect 513 6895 517 6951
rect 453 6891 517 6895
rect 23289 6951 23353 6955
rect 23289 6895 23293 6951
rect 23293 6895 23349 6951
rect 23349 6895 23353 6951
rect 23289 6891 23353 6895
rect 453 6635 517 6639
rect 453 6579 457 6635
rect 457 6579 513 6635
rect 513 6579 517 6635
rect 453 6575 517 6579
rect 23289 6635 23353 6639
rect 23289 6579 23293 6635
rect 23293 6579 23349 6635
rect 23349 6579 23353 6635
rect 23289 6575 23353 6579
rect 453 6398 517 6402
rect 453 6342 457 6398
rect 457 6342 513 6398
rect 513 6342 517 6398
rect 453 6338 517 6342
rect 23289 6398 23353 6402
rect 23289 6342 23293 6398
rect 23293 6342 23349 6398
rect 23349 6342 23353 6398
rect 23289 6338 23353 6342
rect 453 6161 517 6165
rect 453 6105 457 6161
rect 457 6105 513 6161
rect 513 6105 517 6161
rect 453 6101 517 6105
rect 23289 6161 23353 6165
rect 23289 6105 23293 6161
rect 23293 6105 23349 6161
rect 23349 6105 23353 6161
rect 23289 6101 23353 6105
rect 453 5845 517 5849
rect 453 5789 457 5845
rect 457 5789 513 5845
rect 513 5789 517 5845
rect 453 5785 517 5789
rect 23289 5845 23353 5849
rect 23289 5789 23293 5845
rect 23293 5789 23349 5845
rect 23349 5789 23353 5845
rect 23289 5785 23353 5789
rect 453 5608 517 5612
rect 453 5552 457 5608
rect 457 5552 513 5608
rect 513 5552 517 5608
rect 453 5548 517 5552
rect 23289 5608 23353 5612
rect 23289 5552 23293 5608
rect 23293 5552 23349 5608
rect 23349 5552 23353 5608
rect 23289 5548 23353 5552
rect 453 5371 517 5375
rect 453 5315 457 5371
rect 457 5315 513 5371
rect 513 5315 517 5371
rect 453 5311 517 5315
rect 23289 5371 23353 5375
rect 23289 5315 23293 5371
rect 23293 5315 23349 5371
rect 23349 5315 23353 5371
rect 23289 5311 23353 5315
rect 453 5055 517 5059
rect 453 4999 457 5055
rect 457 4999 513 5055
rect 513 4999 517 5055
rect 453 4995 517 4999
rect 23289 5055 23353 5059
rect 23289 4999 23293 5055
rect 23293 4999 23349 5055
rect 23349 4999 23353 5055
rect 23289 4995 23353 4999
rect 453 4818 517 4822
rect 453 4762 457 4818
rect 457 4762 513 4818
rect 513 4762 517 4818
rect 453 4758 517 4762
rect 23289 4818 23353 4822
rect 23289 4762 23293 4818
rect 23293 4762 23349 4818
rect 23349 4762 23353 4818
rect 23289 4758 23353 4762
rect 453 4581 517 4585
rect 453 4525 457 4581
rect 457 4525 513 4581
rect 513 4525 517 4581
rect 453 4521 517 4525
rect 23289 4581 23353 4585
rect 23289 4525 23293 4581
rect 23293 4525 23349 4581
rect 23349 4525 23353 4581
rect 23289 4521 23353 4525
rect 453 4265 517 4269
rect 453 4209 457 4265
rect 457 4209 513 4265
rect 513 4209 517 4265
rect 453 4205 517 4209
rect 23289 4265 23353 4269
rect 23289 4209 23293 4265
rect 23293 4209 23349 4265
rect 23349 4209 23353 4265
rect 23289 4205 23353 4209
rect 453 4028 517 4032
rect 453 3972 457 4028
rect 457 3972 513 4028
rect 513 3972 517 4028
rect 453 3968 517 3972
rect 23289 4028 23353 4032
rect 23289 3972 23293 4028
rect 23293 3972 23349 4028
rect 23349 3972 23353 4028
rect 23289 3968 23353 3972
rect 453 3791 517 3795
rect 453 3735 457 3791
rect 457 3735 513 3791
rect 513 3735 517 3791
rect 453 3731 517 3735
rect 23289 3791 23353 3795
rect 23289 3735 23293 3791
rect 23293 3735 23349 3791
rect 23349 3735 23353 3791
rect 23289 3731 23353 3735
rect 453 3475 517 3479
rect 453 3419 457 3475
rect 457 3419 513 3475
rect 513 3419 517 3475
rect 453 3415 517 3419
rect 23289 3475 23353 3479
rect 23289 3419 23293 3475
rect 23293 3419 23349 3475
rect 23349 3419 23353 3475
rect 23289 3415 23353 3419
rect 453 3238 517 3242
rect 453 3182 457 3238
rect 457 3182 513 3238
rect 513 3182 517 3238
rect 453 3178 517 3182
rect 23289 3238 23353 3242
rect 23289 3182 23293 3238
rect 23293 3182 23349 3238
rect 23349 3182 23353 3238
rect 23289 3178 23353 3182
rect 453 3001 517 3005
rect 453 2945 457 3001
rect 457 2945 513 3001
rect 513 2945 517 3001
rect 453 2941 517 2945
rect 23289 3001 23353 3005
rect 23289 2945 23293 3001
rect 23293 2945 23349 3001
rect 23349 2945 23353 3001
rect 23289 2941 23353 2945
rect 453 2685 517 2689
rect 453 2629 457 2685
rect 457 2629 513 2685
rect 513 2629 517 2685
rect 453 2625 517 2629
rect 23289 2685 23353 2689
rect 23289 2629 23293 2685
rect 23293 2629 23349 2685
rect 23349 2629 23353 2685
rect 23289 2625 23353 2629
rect 453 2448 517 2452
rect 453 2392 457 2448
rect 457 2392 513 2448
rect 513 2392 517 2448
rect 453 2388 517 2392
rect 23289 2448 23353 2452
rect 23289 2392 23293 2448
rect 23293 2392 23349 2448
rect 23349 2392 23353 2448
rect 23289 2388 23353 2392
rect 453 2211 517 2215
rect 453 2155 457 2211
rect 457 2155 513 2211
rect 513 2155 517 2211
rect 453 2151 517 2155
rect 23289 2211 23353 2215
rect 23289 2155 23293 2211
rect 23293 2155 23349 2211
rect 23349 2155 23353 2211
rect 23289 2151 23353 2155
rect 453 1895 517 1899
rect 453 1839 457 1895
rect 457 1839 513 1895
rect 513 1839 517 1895
rect 453 1835 517 1839
rect 23289 1895 23353 1899
rect 23289 1839 23293 1895
rect 23293 1839 23349 1895
rect 23349 1839 23353 1895
rect 23289 1835 23353 1839
rect 453 1658 517 1662
rect 453 1602 457 1658
rect 457 1602 513 1658
rect 513 1602 517 1658
rect 453 1598 517 1602
rect 23289 1658 23353 1662
rect 23289 1602 23293 1658
rect 23293 1602 23349 1658
rect 23349 1602 23353 1658
rect 23289 1598 23353 1602
rect 453 1421 517 1425
rect 453 1365 457 1421
rect 457 1365 513 1421
rect 513 1365 517 1421
rect 453 1361 517 1365
rect 23289 1421 23353 1425
rect 23289 1365 23293 1421
rect 23293 1365 23349 1421
rect 23349 1365 23353 1421
rect 23289 1361 23353 1365
rect 453 1105 517 1109
rect 453 1049 457 1105
rect 457 1049 513 1105
rect 513 1049 517 1105
rect 453 1045 517 1049
rect 23289 1105 23353 1109
rect 23289 1049 23293 1105
rect 23293 1049 23349 1105
rect 23349 1049 23353 1105
rect 23289 1045 23353 1049
rect 453 868 517 872
rect 453 812 457 868
rect 457 812 513 868
rect 513 812 517 868
rect 453 808 517 812
rect 23289 868 23353 872
rect 23289 812 23293 868
rect 23293 812 23349 868
rect 23349 812 23353 868
rect 23289 808 23353 812
rect 453 741 517 745
rect 453 685 457 741
rect 457 685 513 741
rect 513 685 517 741
rect 453 681 517 685
rect 23289 741 23353 745
rect 23289 685 23293 741
rect 23293 685 23349 741
rect 23349 685 23353 741
rect 23289 681 23353 685
rect 43 307 107 311
rect 43 251 47 307
rect 47 251 103 307
rect 103 251 107 307
rect 43 247 107 251
rect 23699 307 23763 311
rect 23699 251 23703 307
rect 23703 251 23759 307
rect 23759 251 23763 307
rect 23699 247 23763 251
<< metal4 >>
rect 42 26713 108 26910
rect 42 26649 43 26713
rect 107 26649 108 26713
rect 42 311 108 26649
rect 42 247 43 311
rect 107 247 108 311
rect 42 0 108 247
rect 452 26499 518 26910
rect 452 26435 453 26499
rect 517 26435 518 26499
rect 452 26152 518 26435
rect 452 26088 453 26152
rect 517 26088 518 26152
rect 452 25915 518 26088
rect 452 25851 453 25915
rect 517 25851 518 25915
rect 452 25599 518 25851
rect 452 25535 453 25599
rect 517 25535 518 25599
rect 452 25362 518 25535
rect 452 25298 453 25362
rect 517 25298 518 25362
rect 452 25125 518 25298
rect 452 25061 453 25125
rect 517 25061 518 25125
rect 452 24809 518 25061
rect 452 24745 453 24809
rect 517 24745 518 24809
rect 452 24572 518 24745
rect 452 24508 453 24572
rect 517 24508 518 24572
rect 452 24335 518 24508
rect 452 24271 453 24335
rect 517 24271 518 24335
rect 452 24019 518 24271
rect 452 23955 453 24019
rect 517 23955 518 24019
rect 452 23782 518 23955
rect 452 23718 453 23782
rect 517 23718 518 23782
rect 452 23545 518 23718
rect 452 23481 453 23545
rect 517 23481 518 23545
rect 452 23229 518 23481
rect 452 23165 453 23229
rect 517 23165 518 23229
rect 452 22992 518 23165
rect 452 22928 453 22992
rect 517 22928 518 22992
rect 452 22755 518 22928
rect 452 22691 453 22755
rect 517 22691 518 22755
rect 452 22439 518 22691
rect 452 22375 453 22439
rect 517 22375 518 22439
rect 452 22202 518 22375
rect 452 22138 453 22202
rect 517 22138 518 22202
rect 452 21965 518 22138
rect 452 21901 453 21965
rect 517 21901 518 21965
rect 452 21649 518 21901
rect 452 21585 453 21649
rect 517 21585 518 21649
rect 452 21412 518 21585
rect 452 21348 453 21412
rect 517 21348 518 21412
rect 452 21175 518 21348
rect 452 21111 453 21175
rect 517 21111 518 21175
rect 452 20859 518 21111
rect 452 20795 453 20859
rect 517 20795 518 20859
rect 452 20622 518 20795
rect 452 20558 453 20622
rect 517 20558 518 20622
rect 452 20385 518 20558
rect 452 20321 453 20385
rect 517 20321 518 20385
rect 452 20069 518 20321
rect 452 20005 453 20069
rect 517 20005 518 20069
rect 452 19832 518 20005
rect 452 19768 453 19832
rect 517 19768 518 19832
rect 452 19595 518 19768
rect 452 19531 453 19595
rect 517 19531 518 19595
rect 452 19279 518 19531
rect 452 19215 453 19279
rect 517 19215 518 19279
rect 452 19042 518 19215
rect 452 18978 453 19042
rect 517 18978 518 19042
rect 452 18805 518 18978
rect 452 18741 453 18805
rect 517 18741 518 18805
rect 452 18489 518 18741
rect 452 18425 453 18489
rect 517 18425 518 18489
rect 452 18252 518 18425
rect 452 18188 453 18252
rect 517 18188 518 18252
rect 452 18015 518 18188
rect 452 17951 453 18015
rect 517 17951 518 18015
rect 452 17699 518 17951
rect 452 17635 453 17699
rect 517 17635 518 17699
rect 452 17462 518 17635
rect 452 17398 453 17462
rect 517 17398 518 17462
rect 452 17225 518 17398
rect 452 17161 453 17225
rect 517 17161 518 17225
rect 452 16909 518 17161
rect 452 16845 453 16909
rect 517 16845 518 16909
rect 452 16672 518 16845
rect 452 16608 453 16672
rect 517 16608 518 16672
rect 452 16435 518 16608
rect 452 16371 453 16435
rect 517 16371 518 16435
rect 452 16119 518 16371
rect 452 16055 453 16119
rect 517 16055 518 16119
rect 452 15882 518 16055
rect 452 15818 453 15882
rect 517 15818 518 15882
rect 452 15645 518 15818
rect 452 15581 453 15645
rect 517 15581 518 15645
rect 452 15329 518 15581
rect 452 15265 453 15329
rect 517 15265 518 15329
rect 452 15092 518 15265
rect 452 15028 453 15092
rect 517 15028 518 15092
rect 452 14855 518 15028
rect 452 14791 453 14855
rect 517 14791 518 14855
rect 452 14539 518 14791
rect 452 14475 453 14539
rect 517 14475 518 14539
rect 452 14302 518 14475
rect 452 14238 453 14302
rect 517 14238 518 14302
rect 452 14065 518 14238
rect 452 14001 453 14065
rect 517 14001 518 14065
rect 452 13749 518 14001
rect 452 13685 453 13749
rect 517 13685 518 13749
rect 452 13512 518 13685
rect 452 13448 453 13512
rect 517 13448 518 13512
rect 452 13275 518 13448
rect 452 13211 453 13275
rect 517 13211 518 13275
rect 452 12959 518 13211
rect 452 12895 453 12959
rect 517 12895 518 12959
rect 452 12722 518 12895
rect 452 12658 453 12722
rect 517 12658 518 12722
rect 452 12485 518 12658
rect 452 12421 453 12485
rect 517 12421 518 12485
rect 452 12169 518 12421
rect 452 12105 453 12169
rect 517 12105 518 12169
rect 452 11932 518 12105
rect 452 11868 453 11932
rect 517 11868 518 11932
rect 452 11695 518 11868
rect 452 11631 453 11695
rect 517 11631 518 11695
rect 452 11379 518 11631
rect 452 11315 453 11379
rect 517 11315 518 11379
rect 452 11142 518 11315
rect 452 11078 453 11142
rect 517 11078 518 11142
rect 452 10905 518 11078
rect 452 10841 453 10905
rect 517 10841 518 10905
rect 452 10589 518 10841
rect 452 10525 453 10589
rect 517 10525 518 10589
rect 452 10352 518 10525
rect 452 10288 453 10352
rect 517 10288 518 10352
rect 452 10115 518 10288
rect 452 10051 453 10115
rect 517 10051 518 10115
rect 452 9799 518 10051
rect 452 9735 453 9799
rect 517 9735 518 9799
rect 452 9562 518 9735
rect 452 9498 453 9562
rect 517 9498 518 9562
rect 452 9325 518 9498
rect 452 9261 453 9325
rect 517 9261 518 9325
rect 452 9009 518 9261
rect 452 8945 453 9009
rect 517 8945 518 9009
rect 452 8772 518 8945
rect 452 8708 453 8772
rect 517 8708 518 8772
rect 452 8535 518 8708
rect 452 8471 453 8535
rect 517 8471 518 8535
rect 452 8219 518 8471
rect 452 8155 453 8219
rect 517 8155 518 8219
rect 452 7982 518 8155
rect 452 7918 453 7982
rect 517 7918 518 7982
rect 452 7745 518 7918
rect 452 7681 453 7745
rect 517 7681 518 7745
rect 452 7429 518 7681
rect 452 7365 453 7429
rect 517 7365 518 7429
rect 452 7192 518 7365
rect 452 7128 453 7192
rect 517 7128 518 7192
rect 452 6955 518 7128
rect 452 6891 453 6955
rect 517 6891 518 6955
rect 452 6639 518 6891
rect 452 6575 453 6639
rect 517 6575 518 6639
rect 452 6402 518 6575
rect 452 6338 453 6402
rect 517 6338 518 6402
rect 452 6165 518 6338
rect 452 6101 453 6165
rect 517 6101 518 6165
rect 452 5849 518 6101
rect 452 5785 453 5849
rect 517 5785 518 5849
rect 452 5612 518 5785
rect 452 5548 453 5612
rect 517 5548 518 5612
rect 452 5375 518 5548
rect 452 5311 453 5375
rect 517 5311 518 5375
rect 452 5059 518 5311
rect 452 4995 453 5059
rect 517 4995 518 5059
rect 452 4822 518 4995
rect 452 4758 453 4822
rect 517 4758 518 4822
rect 452 4585 518 4758
rect 452 4521 453 4585
rect 517 4521 518 4585
rect 452 4269 518 4521
rect 452 4205 453 4269
rect 517 4205 518 4269
rect 452 4032 518 4205
rect 452 3968 453 4032
rect 517 3968 518 4032
rect 452 3795 518 3968
rect 452 3731 453 3795
rect 517 3731 518 3795
rect 452 3479 518 3731
rect 452 3415 453 3479
rect 517 3415 518 3479
rect 452 3242 518 3415
rect 452 3178 453 3242
rect 517 3178 518 3242
rect 452 3005 518 3178
rect 452 2941 453 3005
rect 517 2941 518 3005
rect 452 2689 518 2941
rect 452 2625 453 2689
rect 517 2625 518 2689
rect 452 2452 518 2625
rect 452 2388 453 2452
rect 517 2388 518 2452
rect 452 2215 518 2388
rect 452 2151 453 2215
rect 517 2151 518 2215
rect 452 1899 518 2151
rect 452 1835 453 1899
rect 517 1835 518 1899
rect 452 1662 518 1835
rect 452 1598 453 1662
rect 517 1598 518 1662
rect 452 1425 518 1598
rect 452 1361 453 1425
rect 517 1361 518 1425
rect 452 1109 518 1361
rect 452 1045 453 1109
rect 517 1045 518 1109
rect 452 872 518 1045
rect 452 808 453 872
rect 517 808 518 872
rect 452 745 518 808
rect 452 681 453 745
rect 517 681 518 745
rect 452 0 518 681
rect 23288 26499 23354 26910
rect 23288 26435 23289 26499
rect 23353 26435 23354 26499
rect 23288 26152 23354 26435
rect 23288 26088 23289 26152
rect 23353 26088 23354 26152
rect 23288 25915 23354 26088
rect 23288 25851 23289 25915
rect 23353 25851 23354 25915
rect 23288 25599 23354 25851
rect 23288 25535 23289 25599
rect 23353 25535 23354 25599
rect 23288 25362 23354 25535
rect 23288 25298 23289 25362
rect 23353 25298 23354 25362
rect 23288 25125 23354 25298
rect 23288 25061 23289 25125
rect 23353 25061 23354 25125
rect 23288 24809 23354 25061
rect 23288 24745 23289 24809
rect 23353 24745 23354 24809
rect 23288 24572 23354 24745
rect 23288 24508 23289 24572
rect 23353 24508 23354 24572
rect 23288 24335 23354 24508
rect 23288 24271 23289 24335
rect 23353 24271 23354 24335
rect 23288 24019 23354 24271
rect 23288 23955 23289 24019
rect 23353 23955 23354 24019
rect 23288 23782 23354 23955
rect 23288 23718 23289 23782
rect 23353 23718 23354 23782
rect 23288 23545 23354 23718
rect 23288 23481 23289 23545
rect 23353 23481 23354 23545
rect 23288 23229 23354 23481
rect 23288 23165 23289 23229
rect 23353 23165 23354 23229
rect 23288 22992 23354 23165
rect 23288 22928 23289 22992
rect 23353 22928 23354 22992
rect 23288 22755 23354 22928
rect 23288 22691 23289 22755
rect 23353 22691 23354 22755
rect 23288 22439 23354 22691
rect 23288 22375 23289 22439
rect 23353 22375 23354 22439
rect 23288 22202 23354 22375
rect 23288 22138 23289 22202
rect 23353 22138 23354 22202
rect 23288 21965 23354 22138
rect 23288 21901 23289 21965
rect 23353 21901 23354 21965
rect 23288 21649 23354 21901
rect 23288 21585 23289 21649
rect 23353 21585 23354 21649
rect 23288 21412 23354 21585
rect 23288 21348 23289 21412
rect 23353 21348 23354 21412
rect 23288 21175 23354 21348
rect 23288 21111 23289 21175
rect 23353 21111 23354 21175
rect 23288 20859 23354 21111
rect 23288 20795 23289 20859
rect 23353 20795 23354 20859
rect 23288 20622 23354 20795
rect 23288 20558 23289 20622
rect 23353 20558 23354 20622
rect 23288 20385 23354 20558
rect 23288 20321 23289 20385
rect 23353 20321 23354 20385
rect 23288 20069 23354 20321
rect 23288 20005 23289 20069
rect 23353 20005 23354 20069
rect 23288 19832 23354 20005
rect 23288 19768 23289 19832
rect 23353 19768 23354 19832
rect 23288 19595 23354 19768
rect 23288 19531 23289 19595
rect 23353 19531 23354 19595
rect 23288 19279 23354 19531
rect 23288 19215 23289 19279
rect 23353 19215 23354 19279
rect 23288 19042 23354 19215
rect 23288 18978 23289 19042
rect 23353 18978 23354 19042
rect 23288 18805 23354 18978
rect 23288 18741 23289 18805
rect 23353 18741 23354 18805
rect 23288 18489 23354 18741
rect 23288 18425 23289 18489
rect 23353 18425 23354 18489
rect 23288 18252 23354 18425
rect 23288 18188 23289 18252
rect 23353 18188 23354 18252
rect 23288 18015 23354 18188
rect 23288 17951 23289 18015
rect 23353 17951 23354 18015
rect 23288 17699 23354 17951
rect 23288 17635 23289 17699
rect 23353 17635 23354 17699
rect 23288 17462 23354 17635
rect 23288 17398 23289 17462
rect 23353 17398 23354 17462
rect 23288 17225 23354 17398
rect 23288 17161 23289 17225
rect 23353 17161 23354 17225
rect 23288 16909 23354 17161
rect 23288 16845 23289 16909
rect 23353 16845 23354 16909
rect 23288 16672 23354 16845
rect 23288 16608 23289 16672
rect 23353 16608 23354 16672
rect 23288 16435 23354 16608
rect 23288 16371 23289 16435
rect 23353 16371 23354 16435
rect 23288 16119 23354 16371
rect 23288 16055 23289 16119
rect 23353 16055 23354 16119
rect 23288 15882 23354 16055
rect 23288 15818 23289 15882
rect 23353 15818 23354 15882
rect 23288 15645 23354 15818
rect 23288 15581 23289 15645
rect 23353 15581 23354 15645
rect 23288 15329 23354 15581
rect 23288 15265 23289 15329
rect 23353 15265 23354 15329
rect 23288 15092 23354 15265
rect 23288 15028 23289 15092
rect 23353 15028 23354 15092
rect 23288 14855 23354 15028
rect 23288 14791 23289 14855
rect 23353 14791 23354 14855
rect 23288 14539 23354 14791
rect 23288 14475 23289 14539
rect 23353 14475 23354 14539
rect 23288 14302 23354 14475
rect 23288 14238 23289 14302
rect 23353 14238 23354 14302
rect 23288 14065 23354 14238
rect 23288 14001 23289 14065
rect 23353 14001 23354 14065
rect 23288 13749 23354 14001
rect 23288 13685 23289 13749
rect 23353 13685 23354 13749
rect 23288 13512 23354 13685
rect 23288 13448 23289 13512
rect 23353 13448 23354 13512
rect 23288 13275 23354 13448
rect 23288 13211 23289 13275
rect 23353 13211 23354 13275
rect 23288 12959 23354 13211
rect 23288 12895 23289 12959
rect 23353 12895 23354 12959
rect 23288 12722 23354 12895
rect 23288 12658 23289 12722
rect 23353 12658 23354 12722
rect 23288 12485 23354 12658
rect 23288 12421 23289 12485
rect 23353 12421 23354 12485
rect 23288 12169 23354 12421
rect 23288 12105 23289 12169
rect 23353 12105 23354 12169
rect 23288 11932 23354 12105
rect 23288 11868 23289 11932
rect 23353 11868 23354 11932
rect 23288 11695 23354 11868
rect 23288 11631 23289 11695
rect 23353 11631 23354 11695
rect 23288 11379 23354 11631
rect 23288 11315 23289 11379
rect 23353 11315 23354 11379
rect 23288 11142 23354 11315
rect 23288 11078 23289 11142
rect 23353 11078 23354 11142
rect 23288 10905 23354 11078
rect 23288 10841 23289 10905
rect 23353 10841 23354 10905
rect 23288 10589 23354 10841
rect 23288 10525 23289 10589
rect 23353 10525 23354 10589
rect 23288 10352 23354 10525
rect 23288 10288 23289 10352
rect 23353 10288 23354 10352
rect 23288 10115 23354 10288
rect 23288 10051 23289 10115
rect 23353 10051 23354 10115
rect 23288 9799 23354 10051
rect 23288 9735 23289 9799
rect 23353 9735 23354 9799
rect 23288 9562 23354 9735
rect 23288 9498 23289 9562
rect 23353 9498 23354 9562
rect 23288 9325 23354 9498
rect 23288 9261 23289 9325
rect 23353 9261 23354 9325
rect 23288 9009 23354 9261
rect 23288 8945 23289 9009
rect 23353 8945 23354 9009
rect 23288 8772 23354 8945
rect 23288 8708 23289 8772
rect 23353 8708 23354 8772
rect 23288 8535 23354 8708
rect 23288 8471 23289 8535
rect 23353 8471 23354 8535
rect 23288 8219 23354 8471
rect 23288 8155 23289 8219
rect 23353 8155 23354 8219
rect 23288 7982 23354 8155
rect 23288 7918 23289 7982
rect 23353 7918 23354 7982
rect 23288 7745 23354 7918
rect 23288 7681 23289 7745
rect 23353 7681 23354 7745
rect 23288 7429 23354 7681
rect 23288 7365 23289 7429
rect 23353 7365 23354 7429
rect 23288 7192 23354 7365
rect 23288 7128 23289 7192
rect 23353 7128 23354 7192
rect 23288 6955 23354 7128
rect 23288 6891 23289 6955
rect 23353 6891 23354 6955
rect 23288 6639 23354 6891
rect 23288 6575 23289 6639
rect 23353 6575 23354 6639
rect 23288 6402 23354 6575
rect 23288 6338 23289 6402
rect 23353 6338 23354 6402
rect 23288 6165 23354 6338
rect 23288 6101 23289 6165
rect 23353 6101 23354 6165
rect 23288 5849 23354 6101
rect 23288 5785 23289 5849
rect 23353 5785 23354 5849
rect 23288 5612 23354 5785
rect 23288 5548 23289 5612
rect 23353 5548 23354 5612
rect 23288 5375 23354 5548
rect 23288 5311 23289 5375
rect 23353 5311 23354 5375
rect 23288 5059 23354 5311
rect 23288 4995 23289 5059
rect 23353 4995 23354 5059
rect 23288 4822 23354 4995
rect 23288 4758 23289 4822
rect 23353 4758 23354 4822
rect 23288 4585 23354 4758
rect 23288 4521 23289 4585
rect 23353 4521 23354 4585
rect 23288 4269 23354 4521
rect 23288 4205 23289 4269
rect 23353 4205 23354 4269
rect 23288 4032 23354 4205
rect 23288 3968 23289 4032
rect 23353 3968 23354 4032
rect 23288 3795 23354 3968
rect 23288 3731 23289 3795
rect 23353 3731 23354 3795
rect 23288 3479 23354 3731
rect 23288 3415 23289 3479
rect 23353 3415 23354 3479
rect 23288 3242 23354 3415
rect 23288 3178 23289 3242
rect 23353 3178 23354 3242
rect 23288 3005 23354 3178
rect 23288 2941 23289 3005
rect 23353 2941 23354 3005
rect 23288 2689 23354 2941
rect 23288 2625 23289 2689
rect 23353 2625 23354 2689
rect 23288 2452 23354 2625
rect 23288 2388 23289 2452
rect 23353 2388 23354 2452
rect 23288 2215 23354 2388
rect 23288 2151 23289 2215
rect 23353 2151 23354 2215
rect 23288 1899 23354 2151
rect 23288 1835 23289 1899
rect 23353 1835 23354 1899
rect 23288 1662 23354 1835
rect 23288 1598 23289 1662
rect 23353 1598 23354 1662
rect 23288 1425 23354 1598
rect 23288 1361 23289 1425
rect 23353 1361 23354 1425
rect 23288 1109 23354 1361
rect 23288 1045 23289 1109
rect 23353 1045 23354 1109
rect 23288 872 23354 1045
rect 23288 808 23289 872
rect 23353 808 23354 872
rect 23288 745 23354 808
rect 23288 681 23289 745
rect 23353 681 23354 745
rect 23288 0 23354 681
rect 23698 26713 23764 26910
rect 23698 26649 23699 26713
rect 23763 26649 23764 26713
rect 23698 311 23764 26649
rect 23698 247 23699 311
rect 23763 247 23764 311
rect 23698 0 23764 247
use subbyte2_col_cap_array_0  subbyte2_col_cap_array_0_0
timestamp 1543373569
transform 1 0 1295 0 1 50
box 0 0 21216 474
use subbyte2_col_cap_array  subbyte2_col_cap_array_0
timestamp 1543373569
transform 1 0 1295 0 -1 26910
box 0 0 21216 474
use subbyte2_replica_bitcell_array  subbyte2_replica_bitcell_array_0
timestamp 1543373562
transform 1 0 1295 0 1 445
box -26 -26 21242 26096
use subbyte2_row_cap_array  subbyte2_row_cap_array_0
timestamp 1543373569
transform 1 0 671 0 1 50
box -42 419 624 26441
use subbyte2_row_cap_array_0  subbyte2_row_cap_array_0_0
timestamp 1543373569
transform 1 0 22511 0 1 50
box 0 419 666 26441
<< labels >>
rlabel metal2 s 621 469 23185 517 4 rbl_wl_0_0
port 3 nsew
rlabel metal2 s 621 1163 23185 1211 4 wl_0_0
port 5 nsew
rlabel metal2 s 621 943 23185 991 4 wl_1_0
port 7 nsew
rlabel metal2 s 621 1259 23185 1307 4 wl_0_1
port 9 nsew
rlabel metal2 s 621 1479 23185 1527 4 wl_1_1
port 11 nsew
rlabel metal2 s 621 1953 23185 2001 4 wl_0_2
port 13 nsew
rlabel metal2 s 621 1733 23185 1781 4 wl_1_2
port 15 nsew
rlabel metal2 s 621 2049 23185 2097 4 wl_0_3
port 17 nsew
rlabel metal2 s 621 2269 23185 2317 4 wl_1_3
port 19 nsew
rlabel metal2 s 621 2743 23185 2791 4 wl_0_4
port 21 nsew
rlabel metal2 s 621 2523 23185 2571 4 wl_1_4
port 23 nsew
rlabel metal2 s 621 2839 23185 2887 4 wl_0_5
port 25 nsew
rlabel metal2 s 621 3059 23185 3107 4 wl_1_5
port 27 nsew
rlabel metal2 s 621 3533 23185 3581 4 wl_0_6
port 29 nsew
rlabel metal2 s 621 3313 23185 3361 4 wl_1_6
port 31 nsew
rlabel metal2 s 621 3629 23185 3677 4 wl_0_7
port 33 nsew
rlabel metal2 s 621 3849 23185 3897 4 wl_1_7
port 35 nsew
rlabel metal2 s 621 4323 23185 4371 4 wl_0_8
port 37 nsew
rlabel metal2 s 621 4103 23185 4151 4 wl_1_8
port 39 nsew
rlabel metal2 s 621 4419 23185 4467 4 wl_0_9
port 41 nsew
rlabel metal2 s 621 4639 23185 4687 4 wl_1_9
port 43 nsew
rlabel metal2 s 621 5113 23185 5161 4 wl_0_10
port 45 nsew
rlabel metal2 s 621 4893 23185 4941 4 wl_1_10
port 47 nsew
rlabel metal2 s 621 5209 23185 5257 4 wl_0_11
port 49 nsew
rlabel metal2 s 621 5429 23185 5477 4 wl_1_11
port 51 nsew
rlabel metal2 s 621 5903 23185 5951 4 wl_0_12
port 53 nsew
rlabel metal2 s 621 5683 23185 5731 4 wl_1_12
port 55 nsew
rlabel metal2 s 621 5999 23185 6047 4 wl_0_13
port 57 nsew
rlabel metal2 s 621 6219 23185 6267 4 wl_1_13
port 59 nsew
rlabel metal2 s 621 6693 23185 6741 4 wl_0_14
port 61 nsew
rlabel metal2 s 621 6473 23185 6521 4 wl_1_14
port 63 nsew
rlabel metal2 s 621 6789 23185 6837 4 wl_0_15
port 65 nsew
rlabel metal2 s 621 7009 23185 7057 4 wl_1_15
port 67 nsew
rlabel metal2 s 621 7483 23185 7531 4 wl_0_16
port 69 nsew
rlabel metal2 s 621 7263 23185 7311 4 wl_1_16
port 71 nsew
rlabel metal2 s 621 7579 23185 7627 4 wl_0_17
port 73 nsew
rlabel metal2 s 621 7799 23185 7847 4 wl_1_17
port 75 nsew
rlabel metal2 s 621 8273 23185 8321 4 wl_0_18
port 77 nsew
rlabel metal2 s 621 8053 23185 8101 4 wl_1_18
port 79 nsew
rlabel metal2 s 621 8369 23185 8417 4 wl_0_19
port 81 nsew
rlabel metal2 s 621 8589 23185 8637 4 wl_1_19
port 83 nsew
rlabel metal2 s 621 9063 23185 9111 4 wl_0_20
port 85 nsew
rlabel metal2 s 621 8843 23185 8891 4 wl_1_20
port 87 nsew
rlabel metal2 s 621 9159 23185 9207 4 wl_0_21
port 89 nsew
rlabel metal2 s 621 9379 23185 9427 4 wl_1_21
port 91 nsew
rlabel metal2 s 621 9853 23185 9901 4 wl_0_22
port 93 nsew
rlabel metal2 s 621 9633 23185 9681 4 wl_1_22
port 95 nsew
rlabel metal2 s 621 9949 23185 9997 4 wl_0_23
port 97 nsew
rlabel metal2 s 621 10169 23185 10217 4 wl_1_23
port 99 nsew
rlabel metal2 s 621 10643 23185 10691 4 wl_0_24
port 101 nsew
rlabel metal2 s 621 10423 23185 10471 4 wl_1_24
port 103 nsew
rlabel metal2 s 621 10739 23185 10787 4 wl_0_25
port 105 nsew
rlabel metal2 s 621 10959 23185 11007 4 wl_1_25
port 107 nsew
rlabel metal2 s 621 11433 23185 11481 4 wl_0_26
port 109 nsew
rlabel metal2 s 621 11213 23185 11261 4 wl_1_26
port 111 nsew
rlabel metal2 s 621 11529 23185 11577 4 wl_0_27
port 113 nsew
rlabel metal2 s 621 11749 23185 11797 4 wl_1_27
port 115 nsew
rlabel metal2 s 621 12223 23185 12271 4 wl_0_28
port 117 nsew
rlabel metal2 s 621 12003 23185 12051 4 wl_1_28
port 119 nsew
rlabel metal2 s 621 12319 23185 12367 4 wl_0_29
port 121 nsew
rlabel metal2 s 621 12539 23185 12587 4 wl_1_29
port 123 nsew
rlabel metal2 s 621 13013 23185 13061 4 wl_0_30
port 125 nsew
rlabel metal2 s 621 12793 23185 12841 4 wl_1_30
port 127 nsew
rlabel metal2 s 621 13109 23185 13157 4 wl_0_31
port 129 nsew
rlabel metal2 s 621 13329 23185 13377 4 wl_1_31
port 131 nsew
rlabel metal2 s 621 13803 23185 13851 4 wl_0_32
port 133 nsew
rlabel metal2 s 621 13583 23185 13631 4 wl_1_32
port 135 nsew
rlabel metal2 s 621 13899 23185 13947 4 wl_0_33
port 137 nsew
rlabel metal2 s 621 14119 23185 14167 4 wl_1_33
port 139 nsew
rlabel metal2 s 621 14593 23185 14641 4 wl_0_34
port 141 nsew
rlabel metal2 s 621 14373 23185 14421 4 wl_1_34
port 143 nsew
rlabel metal2 s 621 14689 23185 14737 4 wl_0_35
port 145 nsew
rlabel metal2 s 621 14909 23185 14957 4 wl_1_35
port 147 nsew
rlabel metal2 s 621 15383 23185 15431 4 wl_0_36
port 149 nsew
rlabel metal2 s 621 15163 23185 15211 4 wl_1_36
port 151 nsew
rlabel metal2 s 621 15479 23185 15527 4 wl_0_37
port 153 nsew
rlabel metal2 s 621 15699 23185 15747 4 wl_1_37
port 155 nsew
rlabel metal2 s 621 16173 23185 16221 4 wl_0_38
port 157 nsew
rlabel metal2 s 621 15953 23185 16001 4 wl_1_38
port 159 nsew
rlabel metal2 s 621 16269 23185 16317 4 wl_0_39
port 161 nsew
rlabel metal2 s 621 16489 23185 16537 4 wl_1_39
port 163 nsew
rlabel metal2 s 621 16963 23185 17011 4 wl_0_40
port 165 nsew
rlabel metal2 s 621 16743 23185 16791 4 wl_1_40
port 167 nsew
rlabel metal2 s 621 17059 23185 17107 4 wl_0_41
port 169 nsew
rlabel metal2 s 621 17279 23185 17327 4 wl_1_41
port 171 nsew
rlabel metal2 s 621 17753 23185 17801 4 wl_0_42
port 173 nsew
rlabel metal2 s 621 17533 23185 17581 4 wl_1_42
port 175 nsew
rlabel metal2 s 621 17849 23185 17897 4 wl_0_43
port 177 nsew
rlabel metal2 s 621 18069 23185 18117 4 wl_1_43
port 179 nsew
rlabel metal2 s 621 18543 23185 18591 4 wl_0_44
port 181 nsew
rlabel metal2 s 621 18323 23185 18371 4 wl_1_44
port 183 nsew
rlabel metal2 s 621 18639 23185 18687 4 wl_0_45
port 185 nsew
rlabel metal2 s 621 18859 23185 18907 4 wl_1_45
port 187 nsew
rlabel metal2 s 621 19333 23185 19381 4 wl_0_46
port 189 nsew
rlabel metal2 s 621 19113 23185 19161 4 wl_1_46
port 191 nsew
rlabel metal2 s 621 19429 23185 19477 4 wl_0_47
port 193 nsew
rlabel metal2 s 621 19649 23185 19697 4 wl_1_47
port 195 nsew
rlabel metal2 s 621 20123 23185 20171 4 wl_0_48
port 197 nsew
rlabel metal2 s 621 19903 23185 19951 4 wl_1_48
port 199 nsew
rlabel metal2 s 621 20219 23185 20267 4 wl_0_49
port 201 nsew
rlabel metal2 s 621 20439 23185 20487 4 wl_1_49
port 203 nsew
rlabel metal2 s 621 20913 23185 20961 4 wl_0_50
port 205 nsew
rlabel metal2 s 621 20693 23185 20741 4 wl_1_50
port 207 nsew
rlabel metal2 s 621 21009 23185 21057 4 wl_0_51
port 209 nsew
rlabel metal2 s 621 21229 23185 21277 4 wl_1_51
port 211 nsew
rlabel metal2 s 621 21703 23185 21751 4 wl_0_52
port 213 nsew
rlabel metal2 s 621 21483 23185 21531 4 wl_1_52
port 215 nsew
rlabel metal2 s 621 21799 23185 21847 4 wl_0_53
port 217 nsew
rlabel metal2 s 621 22019 23185 22067 4 wl_1_53
port 219 nsew
rlabel metal2 s 621 22493 23185 22541 4 wl_0_54
port 221 nsew
rlabel metal2 s 621 22273 23185 22321 4 wl_1_54
port 223 nsew
rlabel metal2 s 621 22589 23185 22637 4 wl_0_55
port 225 nsew
rlabel metal2 s 621 22809 23185 22857 4 wl_1_55
port 227 nsew
rlabel metal2 s 621 23283 23185 23331 4 wl_0_56
port 229 nsew
rlabel metal2 s 621 23063 23185 23111 4 wl_1_56
port 231 nsew
rlabel metal2 s 621 23379 23185 23427 4 wl_0_57
port 233 nsew
rlabel metal2 s 621 23599 23185 23647 4 wl_1_57
port 235 nsew
rlabel metal2 s 621 24073 23185 24121 4 wl_0_58
port 237 nsew
rlabel metal2 s 621 23853 23185 23901 4 wl_1_58
port 239 nsew
rlabel metal2 s 621 24169 23185 24217 4 wl_0_59
port 241 nsew
rlabel metal2 s 621 24389 23185 24437 4 wl_1_59
port 243 nsew
rlabel metal2 s 621 24863 23185 24911 4 wl_0_60
port 245 nsew
rlabel metal2 s 621 24643 23185 24691 4 wl_1_60
port 247 nsew
rlabel metal2 s 621 24959 23185 25007 4 wl_0_61
port 249 nsew
rlabel metal2 s 621 25179 23185 25227 4 wl_1_61
port 251 nsew
rlabel metal2 s 621 25653 23185 25701 4 wl_0_62
port 253 nsew
rlabel metal2 s 621 25433 23185 25481 4 wl_1_62
port 255 nsew
rlabel metal2 s 621 25749 23185 25797 4 wl_0_63
port 257 nsew
rlabel metal2 s 621 25969 23185 26017 4 wl_1_63
port 259 nsew
rlabel metal2 s 621 26223 23185 26271 4 rbl_wl_1_1
port 261 nsew
rlabel metal1 s 1805 0 1841 26910 4 rbl_bl_0_0
port 263 nsew
rlabel metal1 s 1589 0 1625 26910 4 rbl_bl_1_0
port 265 nsew
rlabel metal1 s 1733 0 1769 26910 4 rbl_br_0_0
port 267 nsew
rlabel metal1 s 1517 0 1553 26910 4 rbl_br_1_0
port 269 nsew
rlabel metal1 s 1997 0 2033 26910 4 bl_0_0
port 271 nsew
rlabel metal1 s 2213 0 2249 26910 4 bl_1_0
port 273 nsew
rlabel metal1 s 2069 0 2105 26910 4 br_0_0
port 275 nsew
rlabel metal1 s 2285 0 2321 26910 4 br_1_0
port 277 nsew
rlabel metal1 s 3053 0 3089 26910 4 bl_0_1
port 279 nsew
rlabel metal1 s 2837 0 2873 26910 4 bl_1_1
port 281 nsew
rlabel metal1 s 2981 0 3017 26910 4 br_0_1
port 283 nsew
rlabel metal1 s 2765 0 2801 26910 4 br_1_1
port 285 nsew
rlabel metal1 s 3245 0 3281 26910 4 bl_0_2
port 287 nsew
rlabel metal1 s 3461 0 3497 26910 4 bl_1_2
port 289 nsew
rlabel metal1 s 3317 0 3353 26910 4 br_0_2
port 291 nsew
rlabel metal1 s 3533 0 3569 26910 4 br_1_2
port 293 nsew
rlabel metal1 s 4301 0 4337 26910 4 bl_0_3
port 295 nsew
rlabel metal1 s 4085 0 4121 26910 4 bl_1_3
port 297 nsew
rlabel metal1 s 4229 0 4265 26910 4 br_0_3
port 299 nsew
rlabel metal1 s 4013 0 4049 26910 4 br_1_3
port 301 nsew
rlabel metal1 s 4493 0 4529 26910 4 bl_0_4
port 303 nsew
rlabel metal1 s 4709 0 4745 26910 4 bl_1_4
port 305 nsew
rlabel metal1 s 4565 0 4601 26910 4 br_0_4
port 307 nsew
rlabel metal1 s 4781 0 4817 26910 4 br_1_4
port 309 nsew
rlabel metal1 s 5549 0 5585 26910 4 bl_0_5
port 311 nsew
rlabel metal1 s 5333 0 5369 26910 4 bl_1_5
port 313 nsew
rlabel metal1 s 5477 0 5513 26910 4 br_0_5
port 315 nsew
rlabel metal1 s 5261 0 5297 26910 4 br_1_5
port 317 nsew
rlabel metal1 s 5741 0 5777 26910 4 bl_0_6
port 319 nsew
rlabel metal1 s 5957 0 5993 26910 4 bl_1_6
port 321 nsew
rlabel metal1 s 5813 0 5849 26910 4 br_0_6
port 323 nsew
rlabel metal1 s 6029 0 6065 26910 4 br_1_6
port 325 nsew
rlabel metal1 s 6797 0 6833 26910 4 bl_0_7
port 327 nsew
rlabel metal1 s 6581 0 6617 26910 4 bl_1_7
port 329 nsew
rlabel metal1 s 6725 0 6761 26910 4 br_0_7
port 331 nsew
rlabel metal1 s 6509 0 6545 26910 4 br_1_7
port 333 nsew
rlabel metal1 s 6989 0 7025 26910 4 bl_0_8
port 335 nsew
rlabel metal1 s 7205 0 7241 26910 4 bl_1_8
port 337 nsew
rlabel metal1 s 7061 0 7097 26910 4 br_0_8
port 339 nsew
rlabel metal1 s 7277 0 7313 26910 4 br_1_8
port 341 nsew
rlabel metal1 s 8045 0 8081 26910 4 bl_0_9
port 343 nsew
rlabel metal1 s 7829 0 7865 26910 4 bl_1_9
port 345 nsew
rlabel metal1 s 7973 0 8009 26910 4 br_0_9
port 347 nsew
rlabel metal1 s 7757 0 7793 26910 4 br_1_9
port 349 nsew
rlabel metal1 s 8237 0 8273 26910 4 bl_0_10
port 351 nsew
rlabel metal1 s 8453 0 8489 26910 4 bl_1_10
port 353 nsew
rlabel metal1 s 8309 0 8345 26910 4 br_0_10
port 355 nsew
rlabel metal1 s 8525 0 8561 26910 4 br_1_10
port 357 nsew
rlabel metal1 s 9293 0 9329 26910 4 bl_0_11
port 359 nsew
rlabel metal1 s 9077 0 9113 26910 4 bl_1_11
port 361 nsew
rlabel metal1 s 9221 0 9257 26910 4 br_0_11
port 363 nsew
rlabel metal1 s 9005 0 9041 26910 4 br_1_11
port 365 nsew
rlabel metal1 s 9485 0 9521 26910 4 bl_0_12
port 367 nsew
rlabel metal1 s 9701 0 9737 26910 4 bl_1_12
port 369 nsew
rlabel metal1 s 9557 0 9593 26910 4 br_0_12
port 371 nsew
rlabel metal1 s 9773 0 9809 26910 4 br_1_12
port 373 nsew
rlabel metal1 s 10541 0 10577 26910 4 bl_0_13
port 375 nsew
rlabel metal1 s 10325 0 10361 26910 4 bl_1_13
port 377 nsew
rlabel metal1 s 10469 0 10505 26910 4 br_0_13
port 379 nsew
rlabel metal1 s 10253 0 10289 26910 4 br_1_13
port 381 nsew
rlabel metal1 s 10733 0 10769 26910 4 bl_0_14
port 383 nsew
rlabel metal1 s 10949 0 10985 26910 4 bl_1_14
port 385 nsew
rlabel metal1 s 10805 0 10841 26910 4 br_0_14
port 387 nsew
rlabel metal1 s 11021 0 11057 26910 4 br_1_14
port 389 nsew
rlabel metal1 s 11789 0 11825 26910 4 bl_0_15
port 391 nsew
rlabel metal1 s 11573 0 11609 26910 4 bl_1_15
port 393 nsew
rlabel metal1 s 11717 0 11753 26910 4 br_0_15
port 395 nsew
rlabel metal1 s 11501 0 11537 26910 4 br_1_15
port 397 nsew
rlabel metal1 s 11981 0 12017 26910 4 bl_0_16
port 399 nsew
rlabel metal1 s 12197 0 12233 26910 4 bl_1_16
port 401 nsew
rlabel metal1 s 12053 0 12089 26910 4 br_0_16
port 403 nsew
rlabel metal1 s 12269 0 12305 26910 4 br_1_16
port 405 nsew
rlabel metal1 s 13037 0 13073 26910 4 bl_0_17
port 407 nsew
rlabel metal1 s 12821 0 12857 26910 4 bl_1_17
port 409 nsew
rlabel metal1 s 12965 0 13001 26910 4 br_0_17
port 411 nsew
rlabel metal1 s 12749 0 12785 26910 4 br_1_17
port 413 nsew
rlabel metal1 s 13229 0 13265 26910 4 bl_0_18
port 415 nsew
rlabel metal1 s 13445 0 13481 26910 4 bl_1_18
port 417 nsew
rlabel metal1 s 13301 0 13337 26910 4 br_0_18
port 419 nsew
rlabel metal1 s 13517 0 13553 26910 4 br_1_18
port 421 nsew
rlabel metal1 s 14285 0 14321 26910 4 bl_0_19
port 423 nsew
rlabel metal1 s 14069 0 14105 26910 4 bl_1_19
port 425 nsew
rlabel metal1 s 14213 0 14249 26910 4 br_0_19
port 427 nsew
rlabel metal1 s 13997 0 14033 26910 4 br_1_19
port 429 nsew
rlabel metal1 s 14477 0 14513 26910 4 bl_0_20
port 431 nsew
rlabel metal1 s 14693 0 14729 26910 4 bl_1_20
port 433 nsew
rlabel metal1 s 14549 0 14585 26910 4 br_0_20
port 435 nsew
rlabel metal1 s 14765 0 14801 26910 4 br_1_20
port 437 nsew
rlabel metal1 s 15533 0 15569 26910 4 bl_0_21
port 439 nsew
rlabel metal1 s 15317 0 15353 26910 4 bl_1_21
port 441 nsew
rlabel metal1 s 15461 0 15497 26910 4 br_0_21
port 443 nsew
rlabel metal1 s 15245 0 15281 26910 4 br_1_21
port 445 nsew
rlabel metal1 s 15725 0 15761 26910 4 bl_0_22
port 447 nsew
rlabel metal1 s 15941 0 15977 26910 4 bl_1_22
port 449 nsew
rlabel metal1 s 15797 0 15833 26910 4 br_0_22
port 451 nsew
rlabel metal1 s 16013 0 16049 26910 4 br_1_22
port 453 nsew
rlabel metal1 s 16781 0 16817 26910 4 bl_0_23
port 455 nsew
rlabel metal1 s 16565 0 16601 26910 4 bl_1_23
port 457 nsew
rlabel metal1 s 16709 0 16745 26910 4 br_0_23
port 459 nsew
rlabel metal1 s 16493 0 16529 26910 4 br_1_23
port 461 nsew
rlabel metal1 s 16973 0 17009 26910 4 bl_0_24
port 463 nsew
rlabel metal1 s 17189 0 17225 26910 4 bl_1_24
port 465 nsew
rlabel metal1 s 17045 0 17081 26910 4 br_0_24
port 467 nsew
rlabel metal1 s 17261 0 17297 26910 4 br_1_24
port 469 nsew
rlabel metal1 s 18029 0 18065 26910 4 bl_0_25
port 471 nsew
rlabel metal1 s 17813 0 17849 26910 4 bl_1_25
port 473 nsew
rlabel metal1 s 17957 0 17993 26910 4 br_0_25
port 475 nsew
rlabel metal1 s 17741 0 17777 26910 4 br_1_25
port 477 nsew
rlabel metal1 s 18221 0 18257 26910 4 bl_0_26
port 479 nsew
rlabel metal1 s 18437 0 18473 26910 4 bl_1_26
port 481 nsew
rlabel metal1 s 18293 0 18329 26910 4 br_0_26
port 483 nsew
rlabel metal1 s 18509 0 18545 26910 4 br_1_26
port 485 nsew
rlabel metal1 s 19277 0 19313 26910 4 bl_0_27
port 487 nsew
rlabel metal1 s 19061 0 19097 26910 4 bl_1_27
port 489 nsew
rlabel metal1 s 19205 0 19241 26910 4 br_0_27
port 491 nsew
rlabel metal1 s 18989 0 19025 26910 4 br_1_27
port 493 nsew
rlabel metal1 s 19469 0 19505 26910 4 bl_0_28
port 495 nsew
rlabel metal1 s 19685 0 19721 26910 4 bl_1_28
port 497 nsew
rlabel metal1 s 19541 0 19577 26910 4 br_0_28
port 499 nsew
rlabel metal1 s 19757 0 19793 26910 4 br_1_28
port 501 nsew
rlabel metal1 s 20525 0 20561 26910 4 bl_0_29
port 503 nsew
rlabel metal1 s 20309 0 20345 26910 4 bl_1_29
port 505 nsew
rlabel metal1 s 20453 0 20489 26910 4 br_0_29
port 507 nsew
rlabel metal1 s 20237 0 20273 26910 4 br_1_29
port 509 nsew
rlabel metal1 s 20717 0 20753 26910 4 bl_0_30
port 511 nsew
rlabel metal1 s 20933 0 20969 26910 4 bl_1_30
port 513 nsew
rlabel metal1 s 20789 0 20825 26910 4 br_0_30
port 515 nsew
rlabel metal1 s 21005 0 21041 26910 4 br_1_30
port 517 nsew
rlabel metal1 s 21773 0 21809 26910 4 bl_0_31
port 519 nsew
rlabel metal1 s 21557 0 21593 26910 4 bl_1_31
port 521 nsew
rlabel metal1 s 21701 0 21737 26910 4 br_0_31
port 523 nsew
rlabel metal1 s 21485 0 21521 26910 4 br_1_31
port 525 nsew
rlabel metal1 s 21965 0 22001 26910 4 rbl_bl_0_1
port 527 nsew
rlabel metal1 s 22181 0 22217 26910 4 rbl_bl_1_1
port 529 nsew
rlabel metal1 s 22037 0 22073 26910 4 rbl_br_0_1
port 531 nsew
rlabel metal1 s 22253 0 22289 26910 4 rbl_br_1_1
port 533 nsew
rlabel metal4 s 23288 0 23354 26910 4 gnd
port 535 nsew
rlabel metal4 s 452 0 518 26910 4 gnd
port 535 nsew
rlabel metal4 s 23698 0 23764 26910 4 vdd
port 537 nsew
rlabel metal4 s 42 0 108 26910 4 vdd
port 537 nsew
<< properties >>
string FIXED_BBOX 0 0 23806 26910
<< end >>
