
module aes_enc_core (
	clk_clk,
	reset_reset_n,
	q_export_readdata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[63:0]	q_export_readdata;
endmodule
