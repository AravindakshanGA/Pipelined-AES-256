magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect 823 -4467 5671 3504
<< metal1 >>
rect 4347 2186 4353 2238
rect 4405 2186 4411 2238
rect 4223 696 4229 748
rect 4281 696 4287 748
rect 3251 -2116 3257 -2064
rect 3309 -2076 3315 -2064
rect 4347 -2076 4353 -2064
rect 3309 -2104 4353 -2076
rect 3309 -2116 3315 -2104
rect 4347 -2116 4353 -2104
rect 4405 -2116 4411 -2064
rect 2083 -2218 2089 -2166
rect 2141 -2178 2147 -2166
rect 4223 -2178 4229 -2166
rect 2141 -2206 4229 -2178
rect 2141 -2218 2147 -2206
rect 4223 -2218 4229 -2206
rect 4281 -2218 4287 -2166
<< via1 >>
rect 4353 2186 4405 2238
rect 4229 696 4281 748
rect 3257 -2116 3309 -2064
rect 4353 -2116 4405 -2064
rect 2089 -2218 2141 -2166
rect 4229 -2218 4281 -2166
<< metal2 >>
rect 4353 2238 4405 2244
rect 4353 2180 4405 2186
rect 4229 748 4281 754
rect 4229 690 4281 696
rect 3257 -2064 3309 -2058
rect 3257 -2122 3309 -2116
rect 2089 -2166 2141 -2160
rect 2089 -2224 2141 -2218
rect 2101 -3207 2129 -2224
rect 3269 -3207 3297 -2122
rect 4241 -2160 4269 690
rect 4365 -2058 4393 2180
rect 4353 -2064 4405 -2058
rect 4353 -2122 4405 -2116
rect 4229 -2166 4281 -2160
rect 4229 -2224 4281 -2218
<< properties >>
string FIXED_BBOX 2083 -3207 4411 2244
<< end >>
