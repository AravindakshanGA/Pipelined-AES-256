magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1309 -1309 10640 2727
<< locali >>
rect -17 1431 17 1447
rect -17 1381 17 1397
rect 4655 1431 4689 1447
rect 4655 1381 4689 1397
rect 1151 17 1185 33
rect 1151 -33 1185 -17
rect 5823 17 5857 33
rect 5823 -33 5857 -17
<< viali >>
rect -17 1397 17 1431
rect 4655 1397 4689 1431
rect 1151 -17 1185 17
rect 5823 -17 5857 17
<< metal1 >>
rect -32 1388 -26 1440
rect 26 1388 32 1440
rect 4640 1388 4646 1440
rect 4698 1388 4704 1440
rect 1136 -26 1142 26
rect 1194 -26 1200 26
rect 5808 -26 5814 26
rect 5866 -26 5872 26
<< via1 >>
rect -26 1431 26 1440
rect -26 1397 -17 1431
rect -17 1397 17 1431
rect 17 1397 26 1431
rect -26 1388 26 1397
rect 4646 1431 4698 1440
rect 4646 1397 4655 1431
rect 4655 1397 4689 1431
rect 4689 1397 4698 1431
rect 4646 1388 4698 1397
rect 1142 17 1194 26
rect 1142 -17 1151 17
rect 1151 -17 1185 17
rect 1185 -17 1194 17
rect 1142 -26 1194 -17
rect 5814 17 5866 26
rect 5814 -17 5823 17
rect 5823 -17 5857 17
rect 5857 -17 5866 17
rect 5814 -26 5866 -17
<< metal2 >>
rect -28 1442 28 1451
rect 4644 1442 4700 1451
rect -28 1377 28 1386
rect 137 538 203 590
rect 369 345 397 1414
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 1537 345 1565 1414
rect 2250 609 2316 661
rect 2473 538 2539 590
rect 2705 345 2733 1414
rect 3418 609 3484 661
rect 3641 538 3707 590
rect 3873 345 3901 1414
rect 4644 1377 4700 1386
rect 4586 609 4652 661
rect 4809 538 4875 590
rect 5041 345 5069 1414
rect 5754 609 5820 661
rect 5977 538 6043 590
rect 6209 345 6237 1414
rect 6922 609 6988 661
rect 7145 538 7211 590
rect 7377 345 7405 1414
rect 8090 609 8156 661
rect 8313 538 8379 590
rect 8545 345 8573 1414
rect 9258 609 9324 661
rect 368 336 424 345
rect 368 271 424 280
rect 1536 336 1592 345
rect 1536 271 1592 280
rect 2704 336 2760 345
rect 2704 271 2760 280
rect 3872 336 3928 345
rect 3872 271 3928 280
rect 5040 336 5096 345
rect 5040 271 5096 280
rect 6208 336 6264 345
rect 6208 271 6264 280
rect 7376 336 7432 345
rect 7376 271 7432 280
rect 8544 336 8600 345
rect 8544 271 8600 280
rect 369 0 397 271
rect 1140 28 1196 37
rect 1537 0 1565 271
rect 2705 0 2733 271
rect 3873 0 3901 271
rect 5041 0 5069 271
rect 5812 28 5868 37
rect 1140 -37 1196 -28
rect 6209 0 6237 271
rect 7377 0 7405 271
rect 8545 0 8573 271
rect 5812 -37 5868 -28
<< via2 >>
rect -28 1440 28 1442
rect -28 1388 -26 1440
rect -26 1388 26 1440
rect 26 1388 28 1440
rect 4644 1440 4700 1442
rect -28 1386 28 1388
rect 4644 1388 4646 1440
rect 4646 1388 4698 1440
rect 4698 1388 4700 1440
rect 4644 1386 4700 1388
rect 368 280 424 336
rect 1536 280 1592 336
rect 2704 280 2760 336
rect 3872 280 3928 336
rect 5040 280 5096 336
rect 6208 280 6264 336
rect 7376 280 7432 336
rect 8544 280 8600 336
rect 1140 26 1196 28
rect 1140 -26 1142 26
rect 1142 -26 1194 26
rect 1194 -26 1196 26
rect 5812 26 5868 28
rect 1140 -28 1196 -26
rect 5812 -26 5814 26
rect 5814 -26 5866 26
rect 5866 -26 5868 26
rect 5812 -28 5868 -26
<< metal3 >>
rect -49 1442 49 1463
rect -49 1386 -28 1442
rect 28 1386 49 1442
rect -49 1365 49 1386
rect 4623 1442 4721 1463
rect 4623 1386 4644 1442
rect 4700 1386 4721 1442
rect 4623 1365 4721 1386
rect 363 338 429 341
rect 1531 338 1597 341
rect 2699 338 2765 341
rect 3867 338 3933 341
rect 5035 338 5101 341
rect 6203 338 6269 341
rect 7371 338 7437 341
rect 8539 338 8605 341
rect 0 336 9344 338
rect 0 280 368 336
rect 424 280 1536 336
rect 1592 280 2704 336
rect 2760 280 3872 336
rect 3928 280 5040 336
rect 5096 280 6208 336
rect 6264 280 7376 336
rect 7432 280 8544 336
rect 8600 280 9344 336
rect 0 278 9344 280
rect 363 275 429 278
rect 1531 275 1597 278
rect 2699 275 2765 278
rect 3867 275 3933 278
rect 5035 275 5101 278
rect 6203 275 6269 278
rect 7371 275 7437 278
rect 8539 275 8605 278
rect 1119 28 1217 49
rect 1119 -28 1140 28
rect 1196 -28 1217 28
rect 1119 -49 1217 -28
rect 5791 28 5889 49
rect 5791 -28 5812 28
rect 5868 -28 5889 28
rect 5791 -49 5889 -28
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1438349329
transform 1 0 8176 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1438349329
transform 1 0 7008 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1438349329
transform 1 0 5840 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1438349329
transform 1 0 4672 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_4
timestamp 1438349329
transform 1 0 3504 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_5
timestamp 1438349329
transform 1 0 2336 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_6
timestamp 1438349329
transform 1 0 1168 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_7
timestamp 1438349329
transform 1 0 0 0 1 0
box -36 -43 1204 1467
<< labels >>
rlabel metal3 s -49 1365 49 1463 4 vdd
port 3 nsew
rlabel metal3 s 4623 1365 4721 1463 4 vdd
port 3 nsew
rlabel metal3 s 5791 -49 5889 49 4 gnd
port 5 nsew
rlabel metal3 s 1119 -49 1217 49 4 gnd
port 5 nsew
rlabel metal2 s 137 538 203 590 4 din_0
port 7 nsew
rlabel metal2 s 1082 609 1148 661 4 dout_0
port 9 nsew
rlabel metal2 s 1305 538 1371 590 4 din_1
port 11 nsew
rlabel metal2 s 2250 609 2316 661 4 dout_1
port 13 nsew
rlabel metal2 s 2473 538 2539 590 4 din_2
port 15 nsew
rlabel metal2 s 3418 609 3484 661 4 dout_2
port 17 nsew
rlabel metal2 s 3641 538 3707 590 4 din_3
port 19 nsew
rlabel metal2 s 4586 609 4652 661 4 dout_3
port 21 nsew
rlabel metal2 s 4809 538 4875 590 4 din_4
port 23 nsew
rlabel metal2 s 5754 609 5820 661 4 dout_4
port 25 nsew
rlabel metal2 s 5977 538 6043 590 4 din_5
port 27 nsew
rlabel metal2 s 6922 609 6988 661 4 dout_5
port 29 nsew
rlabel metal2 s 7145 538 7211 590 4 din_6
port 31 nsew
rlabel metal2 s 8090 609 8156 661 4 dout_6
port 33 nsew
rlabel metal2 s 8313 538 8379 590 4 din_7
port 35 nsew
rlabel metal2 s 9258 609 9324 661 4 dout_7
port 37 nsew
rlabel metal3 s 0 278 9344 338 4 clk
port 39 nsew
<< properties >>
string FIXED_BBOX 5807 -37 5873 0
<< end >>
