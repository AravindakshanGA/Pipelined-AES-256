magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect 40057 38418 43821 44601
<< metal1 >>
rect 41441 42042 41447 42094
rect 41499 42082 41505 42094
rect 42497 42082 42503 42094
rect 41499 42054 42503 42082
rect 41499 42042 41505 42054
rect 42497 42042 42503 42054
rect 42555 42042 42561 42094
rect 41441 41174 41447 41226
rect 41499 41174 41505 41226
rect 41317 39684 41323 39736
rect 41375 39684 41381 39736
<< via1 >>
rect 41447 42042 41499 42094
rect 42503 42042 42555 42094
rect 41447 41174 41499 41226
rect 41323 39684 41375 39736
<< metal2 >>
rect 41347 41980 41375 43341
rect 42515 42100 42543 43341
rect 41447 42094 41499 42100
rect 41447 42036 41499 42042
rect 42503 42094 42555 42100
rect 42503 42036 42555 42042
rect 41335 41952 41375 41980
rect 41335 39742 41363 41952
rect 41459 41232 41487 42036
rect 41447 41226 41499 41232
rect 41447 41168 41499 41174
rect 41323 39736 41375 39742
rect 41323 39678 41375 39684
<< properties >>
string FIXED_BBOX 41317 39678 42561 43341
<< end >>
