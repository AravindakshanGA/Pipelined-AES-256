magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 3524 2731
<< nwell >>
rect -36 679 2264 1471
<< locali >>
rect 0 1397 2228 1431
rect 64 636 98 702
rect 547 690 817 724
rect 1042 690 1401 724
rect 1719 690 1753 724
rect 196 652 449 686
rect 547 669 581 690
rect 0 -17 2228 17
use subbyte2_pinv  subbyte2_pinv_0
timestamp 1543373571
transform 1 0 368 0 1 0
box -36 -17 404 1471
use subbyte2_pinv  subbyte2_pinv_1
timestamp 1543373571
transform 1 0 0 0 1 0
box -36 -17 404 1471
use subbyte2_pinv_6  subbyte2_pinv_6_0
timestamp 1543373571
transform 1 0 736 0 1 0
box -36 -17 620 1471
use subbyte2_pinv_7  subbyte2_pinv_7_0
timestamp 1543373571
transform 1 0 1320 0 1 0
box -36 -17 944 1471
<< labels >>
rlabel locali s 1736 707 1736 707 4 Z
port 1 nsew
rlabel locali s 81 669 81 669 4 A
port 2 nsew
rlabel locali s 1114 0 1114 0 4 gnd
port 3 nsew
rlabel locali s 1114 1414 1114 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2228 1414
<< end >>
