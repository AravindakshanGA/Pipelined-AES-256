magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 2042 2731
<< locali >>
rect 0 1397 746 1431
rect 330 686 364 1151
rect 330 652 459 686
rect 557 652 591 686
rect 212 485 246 551
rect 112 237 146 303
rect 0 -17 746 17
use subbyte2_pdriver  subbyte2_pdriver_0
timestamp 1543373571
transform 1 0 378 0 1 0
box -36 -17 404 1471
use subbyte2_pnand2  subbyte2_pnand2_0
timestamp 1543373571
transform 1 0 0 0 1 0
box -36 -17 414 1471
<< labels >>
rlabel locali s 574 669 574 669 4 Z
port 1 nsew
rlabel locali s 129 270 129 270 4 A
port 2 nsew
rlabel locali s 229 518 229 518 4 B
port 3 nsew
rlabel locali s 373 0 373 0 4 gnd
port 4 nsew
rlabel locali s 373 1414 373 1414 4 vdd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 746 1414
<< end >>
