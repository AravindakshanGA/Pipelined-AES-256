magic
tech sky130A
magscale 1 2
timestamp 1543373571
<< checkpaint >>
rect -1296 -1277 3544 2731
<< nwell >>
rect -36 679 2284 1471
<< locali >>
rect 0 1397 2248 1431
rect 64 637 98 703
rect 291 690 773 724
rect 1415 690 1449 724
rect 291 670 325 690
rect 0 -17 2248 17
use subbyte2_pinv_9  subbyte2_pinv_9_0
timestamp 1543373571
transform 1 0 0 0 1 0
box -36 -17 728 1471
use subbyte2_pinv_10  subbyte2_pinv_10_0
timestamp 1543373571
transform 1 0 692 0 1 0
box -36 -17 1592 1471
<< labels >>
rlabel locali s 1432 707 1432 707 4 Z
port 1 nsew
rlabel locali s 81 670 81 670 4 A
port 2 nsew
rlabel locali s 1124 0 1124 0 4 gnd
port 3 nsew
rlabel locali s 1124 1414 1124 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2248 1414
<< end >>
