magic
tech sky130A
magscale 1 2
timestamp 1483185662
<< checkpaint >>
rect -1801 -1260 2197 3816
<< nwell >>
rect -541 564 937 1914
<< pwell >>
rect 158 2435 356 2461
rect 158 2291 494 2435
rect 158 2145 356 2291
rect 70 1963 356 2145
rect 72 501 268 522
rect 72 357 424 501
rect 72 340 268 357
<< nmos >>
rect 242 2305 272 2435
rect 154 1989 184 2119
rect 242 1989 272 2119
rect 156 366 186 496
<< pmos >>
rect 154 1624 184 1876
rect 242 1624 272 1876
rect 154 1002 184 1402
rect 346 1002 376 1402
rect 156 602 186 854
<< ndiff >>
rect 184 2420 242 2435
rect 184 2386 196 2420
rect 230 2386 242 2420
rect 184 2352 242 2386
rect 184 2318 196 2352
rect 230 2318 242 2352
rect 184 2305 242 2318
rect 272 2422 330 2435
rect 272 2388 284 2422
rect 318 2388 330 2422
rect 272 2354 330 2388
rect 272 2320 284 2354
rect 318 2320 330 2354
rect 272 2305 330 2320
rect 96 2107 154 2119
rect 96 2073 108 2107
rect 142 2073 154 2107
rect 96 2039 154 2073
rect 96 2005 108 2039
rect 142 2005 154 2039
rect 96 1989 154 2005
rect 184 2107 242 2119
rect 184 2073 196 2107
rect 230 2073 242 2107
rect 184 2039 242 2073
rect 184 2005 196 2039
rect 230 2005 242 2039
rect 184 1989 242 2005
rect 272 2107 330 2119
rect 272 2073 284 2107
rect 318 2073 330 2107
rect 272 2039 330 2073
rect 272 2005 284 2039
rect 318 2005 330 2039
rect 272 1989 330 2005
rect 98 482 156 496
rect 98 448 110 482
rect 144 448 156 482
rect 98 414 156 448
rect 98 380 110 414
rect 144 380 156 414
rect 98 366 156 380
rect 186 482 242 496
rect 186 448 198 482
rect 232 448 242 482
rect 186 414 242 448
rect 186 380 198 414
rect 232 380 242 414
rect 186 366 242 380
<< pdiff >>
rect 100 1835 154 1876
rect 100 1801 108 1835
rect 142 1801 154 1835
rect 100 1767 154 1801
rect 100 1733 108 1767
rect 142 1733 154 1767
rect 100 1699 154 1733
rect 100 1665 108 1699
rect 142 1665 154 1699
rect 100 1624 154 1665
rect 184 1835 242 1876
rect 184 1801 196 1835
rect 230 1801 242 1835
rect 184 1767 242 1801
rect 184 1733 196 1767
rect 230 1733 242 1767
rect 184 1699 242 1733
rect 184 1665 196 1699
rect 230 1665 242 1699
rect 184 1624 242 1665
rect 272 1835 326 1876
rect 272 1801 284 1835
rect 318 1801 326 1835
rect 272 1767 326 1801
rect 272 1733 284 1767
rect 318 1733 326 1767
rect 272 1699 326 1733
rect 272 1665 284 1699
rect 318 1665 326 1699
rect 272 1624 326 1665
rect 100 1389 154 1402
rect 100 1355 108 1389
rect 142 1355 154 1389
rect 100 1321 154 1355
rect 100 1287 108 1321
rect 142 1287 154 1321
rect 100 1253 154 1287
rect 100 1219 108 1253
rect 142 1219 154 1253
rect 100 1185 154 1219
rect 100 1151 108 1185
rect 142 1151 154 1185
rect 100 1117 154 1151
rect 100 1083 108 1117
rect 142 1083 154 1117
rect 100 1049 154 1083
rect 100 1015 108 1049
rect 142 1015 154 1049
rect 100 1002 154 1015
rect 184 1389 238 1402
rect 184 1355 196 1389
rect 230 1355 238 1389
rect 184 1321 238 1355
rect 184 1287 196 1321
rect 230 1287 238 1321
rect 184 1253 238 1287
rect 184 1219 196 1253
rect 230 1219 238 1253
rect 184 1185 238 1219
rect 184 1151 196 1185
rect 230 1151 238 1185
rect 184 1117 238 1151
rect 184 1083 196 1117
rect 230 1083 238 1117
rect 184 1049 238 1083
rect 184 1015 196 1049
rect 230 1015 238 1049
rect 184 1002 238 1015
rect 292 1389 346 1402
rect 292 1355 300 1389
rect 334 1355 346 1389
rect 292 1321 346 1355
rect 292 1287 300 1321
rect 334 1287 346 1321
rect 292 1253 346 1287
rect 292 1219 300 1253
rect 334 1219 346 1253
rect 292 1185 346 1219
rect 292 1151 300 1185
rect 334 1151 346 1185
rect 292 1117 346 1151
rect 292 1083 300 1117
rect 334 1083 346 1117
rect 292 1049 346 1083
rect 292 1015 300 1049
rect 334 1015 346 1049
rect 292 1002 346 1015
rect 376 1389 430 1402
rect 376 1355 388 1389
rect 422 1355 430 1389
rect 376 1321 430 1355
rect 376 1287 388 1321
rect 422 1287 430 1321
rect 376 1253 430 1287
rect 376 1219 388 1253
rect 422 1219 430 1253
rect 376 1185 430 1219
rect 376 1151 388 1185
rect 422 1151 430 1185
rect 376 1117 430 1151
rect 376 1083 388 1117
rect 422 1083 430 1117
rect 376 1049 430 1083
rect 376 1015 388 1049
rect 422 1015 430 1049
rect 376 1002 430 1015
rect 98 813 156 854
rect 98 779 110 813
rect 144 779 156 813
rect 98 745 156 779
rect 98 711 110 745
rect 144 711 156 745
rect 98 677 156 711
rect 98 643 110 677
rect 144 643 156 677
rect 98 602 156 643
rect 186 813 240 854
rect 186 779 198 813
rect 232 779 240 813
rect 186 745 240 779
rect 186 711 198 745
rect 232 711 240 745
rect 186 677 240 711
rect 186 643 198 677
rect 232 643 240 677
rect 186 602 240 643
<< ndiffc >>
rect 196 2386 230 2420
rect 196 2318 230 2352
rect 284 2388 318 2422
rect 284 2320 318 2354
rect 108 2073 142 2107
rect 108 2005 142 2039
rect 196 2073 230 2107
rect 196 2005 230 2039
rect 284 2073 318 2107
rect 284 2005 318 2039
rect 110 448 144 482
rect 110 380 144 414
rect 198 448 232 482
rect 198 380 232 414
<< pdiffc >>
rect 108 1801 142 1835
rect 108 1733 142 1767
rect 108 1665 142 1699
rect 196 1801 230 1835
rect 196 1733 230 1767
rect 196 1665 230 1699
rect 284 1801 318 1835
rect 284 1733 318 1767
rect 284 1665 318 1699
rect 108 1355 142 1389
rect 108 1287 142 1321
rect 108 1219 142 1253
rect 108 1151 142 1185
rect 108 1083 142 1117
rect 108 1015 142 1049
rect 196 1355 230 1389
rect 196 1287 230 1321
rect 196 1219 230 1253
rect 196 1151 230 1185
rect 196 1083 230 1117
rect 196 1015 230 1049
rect 300 1355 334 1389
rect 300 1287 334 1321
rect 300 1219 334 1253
rect 300 1151 334 1185
rect 300 1083 334 1117
rect 300 1015 334 1049
rect 388 1355 422 1389
rect 388 1287 422 1321
rect 388 1219 422 1253
rect 388 1151 422 1185
rect 388 1083 422 1117
rect 388 1015 422 1049
rect 110 779 144 813
rect 110 711 144 745
rect 110 643 144 677
rect 198 779 232 813
rect 198 711 232 745
rect 198 643 232 677
<< psubdiff >>
rect 434 2385 468 2409
rect 434 2317 468 2351
rect 364 451 398 475
rect 364 383 398 417
<< nsubdiff >>
rect 388 1648 422 1676
rect 388 1590 422 1614
<< psubdiffcont >>
rect 434 2351 468 2385
rect 364 417 398 451
<< nsubdiffcont >>
rect 388 1614 422 1648
<< poly >>
rect 240 2520 274 2526
rect 230 2510 284 2520
rect 230 2476 240 2510
rect 274 2476 284 2510
rect 230 2466 284 2476
rect 240 2460 274 2466
rect 242 2435 272 2460
rect 242 2289 272 2305
rect 26 2259 272 2289
rect 26 1448 56 2259
rect 306 2217 372 2227
rect 154 2187 322 2217
rect 154 2119 184 2187
rect 306 2183 322 2187
rect 356 2183 372 2217
rect 306 2173 372 2183
rect 342 2162 372 2173
rect 242 2119 272 2145
rect 342 2128 376 2162
rect 154 1876 184 1989
rect 242 1876 272 1989
rect 345 1976 375 2128
rect 342 1942 376 1976
rect 154 1598 184 1624
rect 242 1556 272 1624
rect 98 1540 272 1556
rect 98 1506 108 1540
rect 142 1526 272 1540
rect 342 1532 372 1942
rect 142 1506 152 1526
rect 98 1496 152 1506
rect 342 1506 474 1532
rect 342 1502 430 1506
rect 108 1490 142 1496
rect 420 1472 430 1502
rect 464 1472 474 1506
rect 420 1458 474 1472
rect 430 1456 474 1458
rect 26 1418 184 1448
rect 154 1402 184 1418
rect 346 1402 376 1428
rect 154 986 184 1002
rect 346 986 376 1002
rect 154 956 376 986
rect 156 898 432 914
rect 156 884 388 898
rect 156 854 186 884
rect 378 864 388 884
rect 422 864 432 898
rect 378 848 432 864
rect 156 496 186 602
rect 156 336 186 366
<< polycont >>
rect 240 2476 274 2510
rect 322 2183 356 2217
rect 108 1506 142 1540
rect 430 1472 464 1506
rect 388 864 422 898
<< locali >>
rect 106 2511 140 2512
rect 140 2477 240 2510
rect 106 2476 240 2477
rect 274 2476 290 2510
rect 196 2420 230 2442
rect 196 2352 230 2386
rect 108 2107 142 2130
rect 108 2039 142 2073
rect 108 1835 142 2005
rect 196 2107 230 2318
rect 284 2422 318 2442
rect 284 2385 318 2388
rect 434 2385 468 2401
rect 284 2354 434 2385
rect 318 2351 434 2354
rect 284 2301 318 2320
rect 196 2039 230 2073
rect 196 1985 230 2005
rect 284 2183 322 2217
rect 356 2183 374 2217
rect 284 2107 318 2183
rect 284 2039 318 2073
rect 108 1767 142 1801
rect 108 1699 142 1733
rect 108 1540 142 1665
rect 196 1835 230 1880
rect 196 1767 230 1801
rect 196 1699 230 1733
rect 196 1586 230 1665
rect 284 1835 318 2005
rect 284 1767 318 1801
rect 284 1699 318 1733
rect 284 1620 318 1665
rect 352 1614 388 1648
rect 422 1614 438 1648
rect 352 1586 386 1614
rect 196 1552 352 1586
rect 108 1389 142 1506
rect 420 1506 474 1522
rect 420 1490 430 1506
rect 388 1472 430 1490
rect 464 1472 474 1506
rect 388 1456 474 1472
rect 108 1321 142 1355
rect 108 1253 142 1287
rect 108 1185 142 1219
rect 108 1117 142 1151
rect 108 1049 142 1083
rect 108 956 142 1015
rect 196 1389 230 1390
rect 196 1321 230 1355
rect 196 1253 230 1287
rect 196 1185 230 1219
rect 196 1117 230 1151
rect 196 1049 230 1083
rect 196 994 230 1015
rect 300 1389 334 1396
rect 300 1321 334 1355
rect 300 1253 334 1287
rect 300 1185 334 1219
rect 300 1117 334 1151
rect 300 1049 334 1083
rect 300 998 334 1015
rect 388 1389 422 1456
rect 388 1321 422 1355
rect 388 1253 422 1287
rect 388 1185 422 1219
rect 388 1117 422 1151
rect 388 1049 422 1083
rect 388 898 422 1015
rect 110 813 144 858
rect 110 745 144 779
rect 110 677 144 711
rect 110 482 144 643
rect 198 813 232 858
rect 388 848 422 864
rect 198 746 232 779
rect 198 745 364 746
rect 232 712 364 745
rect 198 677 232 711
rect 198 598 232 643
rect 110 414 144 448
rect 110 138 144 380
rect 196 482 232 500
rect 196 448 198 482
rect 364 452 398 467
rect 232 451 398 452
rect 232 448 364 451
rect 196 416 364 448
rect 196 414 232 416
rect 196 380 198 414
rect 196 360 232 380
rect 110 95 144 104
<< viali >>
rect 106 2477 140 2511
rect 434 2317 468 2351
rect 352 1552 386 1586
rect 196 1390 230 1424
rect 300 1396 334 1430
rect 364 712 398 746
rect 364 383 398 417
rect 110 104 144 138
<< metal1 >>
rect 94 2511 152 2524
rect 94 2477 106 2511
rect 140 2477 152 2511
rect 94 2464 152 2477
rect 196 1430 230 2556
rect 272 1442 300 2556
rect 428 2351 474 2379
rect 428 2317 434 2351
rect 468 2317 474 2351
rect 428 2305 474 2317
rect 338 1586 400 1602
rect 338 1552 352 1586
rect 386 1552 400 1586
rect 338 1534 400 1552
rect 272 1430 340 1442
rect 184 1424 242 1430
rect 184 1390 196 1424
rect 230 1390 242 1424
rect 184 1384 242 1390
rect 272 1396 300 1430
rect 334 1396 340 1430
rect 272 1384 340 1396
rect 104 138 150 150
rect 104 104 110 138
rect 144 104 150 138
rect 104 0 150 104
rect 196 0 230 1384
rect 272 0 300 1384
rect 358 746 404 768
rect 358 712 364 746
rect 398 712 404 746
rect 358 692 404 712
rect 358 417 404 445
rect 358 383 364 417
rect 398 383 404 417
rect 358 371 404 383
<< labels >>
rlabel metal1 s 104 0 150 150 4 DOUT
port 3 nsew
rlabel metal1 s 196 1430 230 2556 4 BL
port 5 nsew
rlabel metal1 s 272 1442 300 2556 4 BR
port 7 nsew
rlabel metal1 s 94 2464 152 2524 4 EN
port 9 nsew
rlabel metal1 s 428 2305 474 2379 4 GND
port 11 nsew
rlabel metal1 s 358 371 404 445 4 GND
port 11 nsew
rlabel metal1 s 338 1534 400 1602 4 VDD
port 13 nsew
rlabel metal1 s 358 692 404 768 4 VDD
port 13 nsew
rlabel metal1 s 213 1993 213 1993 4 bl
port 14 nsew
rlabel metal1 s 286 1999 286 1999 4 br
port 15 nsew
rlabel metal1 s 127 75 127 75 4 dout
port 16 nsew
rlabel metal1 s 123 2494 123 2494 4 en
port 17 nsew
rlabel metal1 s 369 1568 369 1568 4 vdd
port 18 nsew
rlabel metal1 s 381 730 381 730 4 vdd
port 18 nsew
rlabel metal1 s 451 2342 451 2342 4 gnd
port 19 nsew
rlabel metal1 s 381 408 381 408 4 gnd
port 19 nsew
<< properties >>
string FIXED_BBOX 0 0 500 2556
<< end >>
