magic
tech sky130A
magscale 1 2
timestamp 1543373570
<< checkpaint >>
rect -1227 -1272 23180 1982
<< locali >>
rect 1709 645 1743 661
rect 1709 595 1743 611
rect 2095 645 2129 661
rect 2095 595 2129 611
rect 2957 645 2991 661
rect 2957 595 2991 611
rect 3343 645 3377 661
rect 3343 595 3377 611
rect 4205 645 4239 661
rect 4205 595 4239 611
rect 4591 645 4625 661
rect 4591 595 4625 611
rect 5453 645 5487 661
rect 5453 595 5487 611
rect 5839 645 5873 661
rect 5839 595 5873 611
rect 6701 645 6735 661
rect 6701 595 6735 611
rect 7087 645 7121 661
rect 7087 595 7121 611
rect 7949 645 7983 661
rect 7949 595 7983 611
rect 8335 645 8369 661
rect 8335 595 8369 611
rect 9197 645 9231 661
rect 9197 595 9231 611
rect 9583 645 9617 661
rect 9583 595 9617 611
rect 10445 645 10479 661
rect 10445 595 10479 611
rect 10831 645 10865 661
rect 10831 595 10865 611
rect 11693 645 11727 661
rect 11693 595 11727 611
rect 12079 645 12113 661
rect 12079 595 12113 611
rect 12941 645 12975 661
rect 12941 595 12975 611
rect 13327 645 13361 661
rect 13327 595 13361 611
rect 14189 645 14223 661
rect 14189 595 14223 611
rect 14575 645 14609 661
rect 14575 595 14609 611
rect 15437 645 15471 661
rect 15437 595 15471 611
rect 15823 645 15857 661
rect 15823 595 15857 611
rect 16685 645 16719 661
rect 16685 595 16719 611
rect 17071 645 17105 661
rect 17071 595 17105 611
rect 17933 645 17967 661
rect 17933 595 17967 611
rect 18319 645 18353 661
rect 18319 595 18353 611
rect 19181 645 19215 661
rect 19181 595 19215 611
rect 19567 645 19601 661
rect 19567 595 19601 611
rect 20429 645 20463 661
rect 20429 595 20463 611
rect 20815 645 20849 661
rect 20815 595 20849 611
rect 21677 645 21711 661
rect 21677 595 21711 611
<< viali >>
rect 1709 611 1743 645
rect 2095 611 2129 645
rect 2957 611 2991 645
rect 3343 611 3377 645
rect 4205 611 4239 645
rect 4591 611 4625 645
rect 5453 611 5487 645
rect 5839 611 5873 645
rect 6701 611 6735 645
rect 7087 611 7121 645
rect 7949 611 7983 645
rect 8335 611 8369 645
rect 9197 611 9231 645
rect 9583 611 9617 645
rect 10445 611 10479 645
rect 10831 611 10865 645
rect 11693 611 11727 645
rect 12079 611 12113 645
rect 12941 611 12975 645
rect 13327 611 13361 645
rect 14189 611 14223 645
rect 14575 611 14609 645
rect 15437 611 15471 645
rect 15823 611 15857 645
rect 16685 611 16719 645
rect 17071 611 17105 645
rect 17933 611 17967 645
rect 18319 611 18353 645
rect 19181 611 19215 645
rect 19567 611 19601 645
rect 20429 611 20463 645
rect 20815 611 20849 645
rect 21677 611 21711 645
<< metal1 >>
rect 1361 0 1389 722
rect 1694 602 1700 654
rect 1752 602 1758 654
rect 1825 0 1853 722
rect 1985 0 2013 722
rect 2080 602 2086 654
rect 2138 602 2144 654
rect 2449 0 2477 722
rect 2609 0 2637 722
rect 2942 602 2948 654
rect 3000 602 3006 654
rect 3073 0 3101 722
rect 3233 0 3261 722
rect 3328 602 3334 654
rect 3386 602 3392 654
rect 3697 0 3725 722
rect 3857 0 3885 722
rect 4190 602 4196 654
rect 4248 602 4254 654
rect 4321 0 4349 722
rect 4481 0 4509 722
rect 4576 602 4582 654
rect 4634 602 4640 654
rect 4945 0 4973 722
rect 5105 0 5133 722
rect 5438 602 5444 654
rect 5496 602 5502 654
rect 5569 0 5597 722
rect 5729 0 5757 722
rect 5824 602 5830 654
rect 5882 602 5888 654
rect 6193 0 6221 722
rect 6353 0 6381 722
rect 6686 602 6692 654
rect 6744 602 6750 654
rect 6817 0 6845 722
rect 6977 0 7005 722
rect 7072 602 7078 654
rect 7130 602 7136 654
rect 7441 0 7469 722
rect 7601 0 7629 722
rect 7934 602 7940 654
rect 7992 602 7998 654
rect 8065 0 8093 722
rect 8225 0 8253 722
rect 8320 602 8326 654
rect 8378 602 8384 654
rect 8689 0 8717 722
rect 8849 0 8877 722
rect 9182 602 9188 654
rect 9240 602 9246 654
rect 9313 0 9341 722
rect 9473 0 9501 722
rect 9568 602 9574 654
rect 9626 602 9632 654
rect 9937 0 9965 722
rect 10097 0 10125 722
rect 10430 602 10436 654
rect 10488 602 10494 654
rect 10561 0 10589 722
rect 10721 0 10749 722
rect 10816 602 10822 654
rect 10874 602 10880 654
rect 11185 0 11213 722
rect 11345 0 11373 722
rect 11678 602 11684 654
rect 11736 602 11742 654
rect 11809 0 11837 722
rect 11969 0 11997 722
rect 12064 602 12070 654
rect 12122 602 12128 654
rect 12433 0 12461 722
rect 12593 0 12621 722
rect 12926 602 12932 654
rect 12984 602 12990 654
rect 13057 0 13085 722
rect 13217 0 13245 722
rect 13312 602 13318 654
rect 13370 602 13376 654
rect 13681 0 13709 722
rect 13841 0 13869 722
rect 14174 602 14180 654
rect 14232 602 14238 654
rect 14305 0 14333 722
rect 14465 0 14493 722
rect 14560 602 14566 654
rect 14618 602 14624 654
rect 14929 0 14957 722
rect 15089 0 15117 722
rect 15422 602 15428 654
rect 15480 602 15486 654
rect 15553 0 15581 722
rect 15713 0 15741 722
rect 15808 602 15814 654
rect 15866 602 15872 654
rect 16177 0 16205 722
rect 16337 0 16365 722
rect 16670 602 16676 654
rect 16728 602 16734 654
rect 16801 0 16829 722
rect 16961 0 16989 722
rect 17056 602 17062 654
rect 17114 602 17120 654
rect 17425 0 17453 722
rect 17585 0 17613 722
rect 17918 602 17924 654
rect 17976 602 17982 654
rect 18049 0 18077 722
rect 18209 0 18237 722
rect 18304 602 18310 654
rect 18362 602 18368 654
rect 18673 0 18701 722
rect 18833 0 18861 722
rect 19166 602 19172 654
rect 19224 602 19230 654
rect 19297 0 19325 722
rect 19457 0 19485 722
rect 19552 602 19558 654
rect 19610 602 19616 654
rect 19921 0 19949 722
rect 20081 0 20109 722
rect 20414 602 20420 654
rect 20472 602 20478 654
rect 20545 0 20573 722
rect 20705 0 20733 722
rect 20800 602 20806 654
rect 20858 602 20864 654
rect 21169 0 21197 722
rect 21329 0 21357 722
rect 21662 602 21668 654
rect 21720 602 21726 654
rect 21793 0 21821 722
<< via1 >>
rect 1700 645 1752 654
rect 1700 611 1709 645
rect 1709 611 1743 645
rect 1743 611 1752 645
rect 1700 602 1752 611
rect 2086 645 2138 654
rect 2086 611 2095 645
rect 2095 611 2129 645
rect 2129 611 2138 645
rect 2086 602 2138 611
rect 2948 645 3000 654
rect 2948 611 2957 645
rect 2957 611 2991 645
rect 2991 611 3000 645
rect 2948 602 3000 611
rect 3334 645 3386 654
rect 3334 611 3343 645
rect 3343 611 3377 645
rect 3377 611 3386 645
rect 3334 602 3386 611
rect 4196 645 4248 654
rect 4196 611 4205 645
rect 4205 611 4239 645
rect 4239 611 4248 645
rect 4196 602 4248 611
rect 4582 645 4634 654
rect 4582 611 4591 645
rect 4591 611 4625 645
rect 4625 611 4634 645
rect 4582 602 4634 611
rect 5444 645 5496 654
rect 5444 611 5453 645
rect 5453 611 5487 645
rect 5487 611 5496 645
rect 5444 602 5496 611
rect 5830 645 5882 654
rect 5830 611 5839 645
rect 5839 611 5873 645
rect 5873 611 5882 645
rect 5830 602 5882 611
rect 6692 645 6744 654
rect 6692 611 6701 645
rect 6701 611 6735 645
rect 6735 611 6744 645
rect 6692 602 6744 611
rect 7078 645 7130 654
rect 7078 611 7087 645
rect 7087 611 7121 645
rect 7121 611 7130 645
rect 7078 602 7130 611
rect 7940 645 7992 654
rect 7940 611 7949 645
rect 7949 611 7983 645
rect 7983 611 7992 645
rect 7940 602 7992 611
rect 8326 645 8378 654
rect 8326 611 8335 645
rect 8335 611 8369 645
rect 8369 611 8378 645
rect 8326 602 8378 611
rect 9188 645 9240 654
rect 9188 611 9197 645
rect 9197 611 9231 645
rect 9231 611 9240 645
rect 9188 602 9240 611
rect 9574 645 9626 654
rect 9574 611 9583 645
rect 9583 611 9617 645
rect 9617 611 9626 645
rect 9574 602 9626 611
rect 10436 645 10488 654
rect 10436 611 10445 645
rect 10445 611 10479 645
rect 10479 611 10488 645
rect 10436 602 10488 611
rect 10822 645 10874 654
rect 10822 611 10831 645
rect 10831 611 10865 645
rect 10865 611 10874 645
rect 10822 602 10874 611
rect 11684 645 11736 654
rect 11684 611 11693 645
rect 11693 611 11727 645
rect 11727 611 11736 645
rect 11684 602 11736 611
rect 12070 645 12122 654
rect 12070 611 12079 645
rect 12079 611 12113 645
rect 12113 611 12122 645
rect 12070 602 12122 611
rect 12932 645 12984 654
rect 12932 611 12941 645
rect 12941 611 12975 645
rect 12975 611 12984 645
rect 12932 602 12984 611
rect 13318 645 13370 654
rect 13318 611 13327 645
rect 13327 611 13361 645
rect 13361 611 13370 645
rect 13318 602 13370 611
rect 14180 645 14232 654
rect 14180 611 14189 645
rect 14189 611 14223 645
rect 14223 611 14232 645
rect 14180 602 14232 611
rect 14566 645 14618 654
rect 14566 611 14575 645
rect 14575 611 14609 645
rect 14609 611 14618 645
rect 14566 602 14618 611
rect 15428 645 15480 654
rect 15428 611 15437 645
rect 15437 611 15471 645
rect 15471 611 15480 645
rect 15428 602 15480 611
rect 15814 645 15866 654
rect 15814 611 15823 645
rect 15823 611 15857 645
rect 15857 611 15866 645
rect 15814 602 15866 611
rect 16676 645 16728 654
rect 16676 611 16685 645
rect 16685 611 16719 645
rect 16719 611 16728 645
rect 16676 602 16728 611
rect 17062 645 17114 654
rect 17062 611 17071 645
rect 17071 611 17105 645
rect 17105 611 17114 645
rect 17062 602 17114 611
rect 17924 645 17976 654
rect 17924 611 17933 645
rect 17933 611 17967 645
rect 17967 611 17976 645
rect 17924 602 17976 611
rect 18310 645 18362 654
rect 18310 611 18319 645
rect 18319 611 18353 645
rect 18353 611 18362 645
rect 18310 602 18362 611
rect 19172 645 19224 654
rect 19172 611 19181 645
rect 19181 611 19215 645
rect 19215 611 19224 645
rect 19172 602 19224 611
rect 19558 645 19610 654
rect 19558 611 19567 645
rect 19567 611 19601 645
rect 19601 611 19610 645
rect 19558 602 19610 611
rect 20420 645 20472 654
rect 20420 611 20429 645
rect 20429 611 20463 645
rect 20463 611 20472 645
rect 20420 602 20472 611
rect 20806 645 20858 654
rect 20806 611 20815 645
rect 20815 611 20849 645
rect 20849 611 20858 645
rect 20806 602 20858 611
rect 21668 645 21720 654
rect 21668 611 21677 645
rect 21677 611 21711 645
rect 21711 611 21720 645
rect 21668 602 21720 611
<< metal2 >>
rect 1698 656 1754 665
rect 1698 591 1754 600
rect 2084 656 2140 665
rect 2084 591 2140 600
rect 2946 656 3002 665
rect 2946 591 3002 600
rect 3332 656 3388 665
rect 3332 591 3388 600
rect 4194 656 4250 665
rect 4194 591 4250 600
rect 4580 656 4636 665
rect 4580 591 4636 600
rect 5442 656 5498 665
rect 5442 591 5498 600
rect 5828 656 5884 665
rect 5828 591 5884 600
rect 6690 656 6746 665
rect 6690 591 6746 600
rect 7076 656 7132 665
rect 7076 591 7132 600
rect 7938 656 7994 665
rect 7938 591 7994 600
rect 8324 656 8380 665
rect 8324 591 8380 600
rect 9186 656 9242 665
rect 9186 591 9242 600
rect 9572 656 9628 665
rect 9572 591 9628 600
rect 10434 656 10490 665
rect 10434 591 10490 600
rect 10820 656 10876 665
rect 10820 591 10876 600
rect 11682 656 11738 665
rect 11682 591 11738 600
rect 12068 656 12124 665
rect 12068 591 12124 600
rect 12930 656 12986 665
rect 12930 591 12986 600
rect 13316 656 13372 665
rect 13316 591 13372 600
rect 14178 656 14234 665
rect 14178 591 14234 600
rect 14564 656 14620 665
rect 14564 591 14620 600
rect 15426 656 15482 665
rect 15426 591 15482 600
rect 15812 656 15868 665
rect 15812 591 15868 600
rect 16674 656 16730 665
rect 16674 591 16730 600
rect 17060 656 17116 665
rect 17060 591 17116 600
rect 17922 656 17978 665
rect 17922 591 17978 600
rect 18308 656 18364 665
rect 18308 591 18364 600
rect 19170 656 19226 665
rect 19170 591 19226 600
rect 19556 656 19612 665
rect 19556 591 19612 600
rect 20418 656 20474 665
rect 20418 591 20474 600
rect 20804 656 20860 665
rect 20804 591 20860 600
rect 21666 656 21722 665
rect 21666 591 21722 600
rect 1579 53 1635 62
rect 1579 -12 1635 -3
rect 2203 53 2259 62
rect 2203 -12 2259 -3
rect 2827 53 2883 62
rect 2827 -12 2883 -3
rect 3451 53 3507 62
rect 3451 -12 3507 -3
rect 4075 53 4131 62
rect 4075 -12 4131 -3
rect 4699 53 4755 62
rect 4699 -12 4755 -3
rect 5323 53 5379 62
rect 5323 -12 5379 -3
rect 5947 53 6003 62
rect 5947 -12 6003 -3
rect 6571 53 6627 62
rect 6571 -12 6627 -3
rect 7195 53 7251 62
rect 7195 -12 7251 -3
rect 7819 53 7875 62
rect 7819 -12 7875 -3
rect 8443 53 8499 62
rect 8443 -12 8499 -3
rect 9067 53 9123 62
rect 9067 -12 9123 -3
rect 9691 53 9747 62
rect 9691 -12 9747 -3
rect 10315 53 10371 62
rect 10315 -12 10371 -3
rect 10939 53 10995 62
rect 10939 -12 10995 -3
rect 11563 53 11619 62
rect 11563 -12 11619 -3
rect 12187 53 12243 62
rect 12187 -12 12243 -3
rect 12811 53 12867 62
rect 12811 -12 12867 -3
rect 13435 53 13491 62
rect 13435 -12 13491 -3
rect 14059 53 14115 62
rect 14059 -12 14115 -3
rect 14683 53 14739 62
rect 14683 -12 14739 -3
rect 15307 53 15363 62
rect 15307 -12 15363 -3
rect 15931 53 15987 62
rect 15931 -12 15987 -3
rect 16555 53 16611 62
rect 16555 -12 16611 -3
rect 17179 53 17235 62
rect 17179 -12 17235 -3
rect 17803 53 17859 62
rect 17803 -12 17859 -3
rect 18427 53 18483 62
rect 18427 -12 18483 -3
rect 19051 53 19107 62
rect 19051 -12 19107 -3
rect 19675 53 19731 62
rect 19675 -12 19731 -3
rect 20299 53 20355 62
rect 20299 -12 20355 -3
rect 20923 53 20979 62
rect 20923 -12 20979 -3
rect 21547 53 21603 62
rect 21547 -12 21603 -3
<< via2 >>
rect 1698 654 1754 656
rect 1698 602 1700 654
rect 1700 602 1752 654
rect 1752 602 1754 654
rect 1698 600 1754 602
rect 2084 654 2140 656
rect 2084 602 2086 654
rect 2086 602 2138 654
rect 2138 602 2140 654
rect 2084 600 2140 602
rect 2946 654 3002 656
rect 2946 602 2948 654
rect 2948 602 3000 654
rect 3000 602 3002 654
rect 2946 600 3002 602
rect 3332 654 3388 656
rect 3332 602 3334 654
rect 3334 602 3386 654
rect 3386 602 3388 654
rect 3332 600 3388 602
rect 4194 654 4250 656
rect 4194 602 4196 654
rect 4196 602 4248 654
rect 4248 602 4250 654
rect 4194 600 4250 602
rect 4580 654 4636 656
rect 4580 602 4582 654
rect 4582 602 4634 654
rect 4634 602 4636 654
rect 4580 600 4636 602
rect 5442 654 5498 656
rect 5442 602 5444 654
rect 5444 602 5496 654
rect 5496 602 5498 654
rect 5442 600 5498 602
rect 5828 654 5884 656
rect 5828 602 5830 654
rect 5830 602 5882 654
rect 5882 602 5884 654
rect 5828 600 5884 602
rect 6690 654 6746 656
rect 6690 602 6692 654
rect 6692 602 6744 654
rect 6744 602 6746 654
rect 6690 600 6746 602
rect 7076 654 7132 656
rect 7076 602 7078 654
rect 7078 602 7130 654
rect 7130 602 7132 654
rect 7076 600 7132 602
rect 7938 654 7994 656
rect 7938 602 7940 654
rect 7940 602 7992 654
rect 7992 602 7994 654
rect 7938 600 7994 602
rect 8324 654 8380 656
rect 8324 602 8326 654
rect 8326 602 8378 654
rect 8378 602 8380 654
rect 8324 600 8380 602
rect 9186 654 9242 656
rect 9186 602 9188 654
rect 9188 602 9240 654
rect 9240 602 9242 654
rect 9186 600 9242 602
rect 9572 654 9628 656
rect 9572 602 9574 654
rect 9574 602 9626 654
rect 9626 602 9628 654
rect 9572 600 9628 602
rect 10434 654 10490 656
rect 10434 602 10436 654
rect 10436 602 10488 654
rect 10488 602 10490 654
rect 10434 600 10490 602
rect 10820 654 10876 656
rect 10820 602 10822 654
rect 10822 602 10874 654
rect 10874 602 10876 654
rect 10820 600 10876 602
rect 11682 654 11738 656
rect 11682 602 11684 654
rect 11684 602 11736 654
rect 11736 602 11738 654
rect 11682 600 11738 602
rect 12068 654 12124 656
rect 12068 602 12070 654
rect 12070 602 12122 654
rect 12122 602 12124 654
rect 12068 600 12124 602
rect 12930 654 12986 656
rect 12930 602 12932 654
rect 12932 602 12984 654
rect 12984 602 12986 654
rect 12930 600 12986 602
rect 13316 654 13372 656
rect 13316 602 13318 654
rect 13318 602 13370 654
rect 13370 602 13372 654
rect 13316 600 13372 602
rect 14178 654 14234 656
rect 14178 602 14180 654
rect 14180 602 14232 654
rect 14232 602 14234 654
rect 14178 600 14234 602
rect 14564 654 14620 656
rect 14564 602 14566 654
rect 14566 602 14618 654
rect 14618 602 14620 654
rect 14564 600 14620 602
rect 15426 654 15482 656
rect 15426 602 15428 654
rect 15428 602 15480 654
rect 15480 602 15482 654
rect 15426 600 15482 602
rect 15812 654 15868 656
rect 15812 602 15814 654
rect 15814 602 15866 654
rect 15866 602 15868 654
rect 15812 600 15868 602
rect 16674 654 16730 656
rect 16674 602 16676 654
rect 16676 602 16728 654
rect 16728 602 16730 654
rect 16674 600 16730 602
rect 17060 654 17116 656
rect 17060 602 17062 654
rect 17062 602 17114 654
rect 17114 602 17116 654
rect 17060 600 17116 602
rect 17922 654 17978 656
rect 17922 602 17924 654
rect 17924 602 17976 654
rect 17976 602 17978 654
rect 17922 600 17978 602
rect 18308 654 18364 656
rect 18308 602 18310 654
rect 18310 602 18362 654
rect 18362 602 18364 654
rect 18308 600 18364 602
rect 19170 654 19226 656
rect 19170 602 19172 654
rect 19172 602 19224 654
rect 19224 602 19226 654
rect 19170 600 19226 602
rect 19556 654 19612 656
rect 19556 602 19558 654
rect 19558 602 19610 654
rect 19610 602 19612 654
rect 19556 600 19612 602
rect 20418 654 20474 656
rect 20418 602 20420 654
rect 20420 602 20472 654
rect 20472 602 20474 654
rect 20418 600 20474 602
rect 20804 654 20860 656
rect 20804 602 20806 654
rect 20806 602 20858 654
rect 20858 602 20860 654
rect 20804 600 20860 602
rect 21666 654 21722 656
rect 21666 602 21668 654
rect 21668 602 21720 654
rect 21720 602 21722 654
rect 21666 600 21722 602
rect 1579 -3 1635 53
rect 2203 -3 2259 53
rect 2827 -3 2883 53
rect 3451 -3 3507 53
rect 4075 -3 4131 53
rect 4699 -3 4755 53
rect 5323 -3 5379 53
rect 5947 -3 6003 53
rect 6571 -3 6627 53
rect 7195 -3 7251 53
rect 7819 -3 7875 53
rect 8443 -3 8499 53
rect 9067 -3 9123 53
rect 9691 -3 9747 53
rect 10315 -3 10371 53
rect 10939 -3 10995 53
rect 11563 -3 11619 53
rect 12187 -3 12243 53
rect 12811 -3 12867 53
rect 13435 -3 13491 53
rect 14059 -3 14115 53
rect 14683 -3 14739 53
rect 15307 -3 15363 53
rect 15931 -3 15987 53
rect 16555 -3 16611 53
rect 17179 -3 17235 53
rect 17803 -3 17859 53
rect 18427 -3 18483 53
rect 19051 -3 19107 53
rect 19675 -3 19731 53
rect 20299 -3 20355 53
rect 20923 -3 20979 53
rect 21547 -3 21603 53
<< metal3 >>
rect 33 656 21920 661
rect 33 600 1698 656
rect 1754 600 2084 656
rect 2140 600 2946 656
rect 3002 600 3332 656
rect 3388 600 4194 656
rect 4250 600 4580 656
rect 4636 600 5442 656
rect 5498 600 5828 656
rect 5884 600 6690 656
rect 6746 600 7076 656
rect 7132 600 7938 656
rect 7994 600 8324 656
rect 8380 600 9186 656
rect 9242 600 9572 656
rect 9628 600 10434 656
rect 10490 600 10820 656
rect 10876 600 11682 656
rect 11738 600 12068 656
rect 12124 600 12930 656
rect 12986 600 13316 656
rect 13372 600 14178 656
rect 14234 600 14564 656
rect 14620 600 15426 656
rect 15482 600 15812 656
rect 15868 600 16674 656
rect 16730 600 17060 656
rect 17116 600 17922 656
rect 17978 600 18308 656
rect 18364 600 19170 656
rect 19226 600 19556 656
rect 19612 600 20418 656
rect 20474 600 20804 656
rect 20860 600 21666 656
rect 21722 600 21920 656
rect 33 595 21920 600
rect 33 53 21920 58
rect 33 -3 1579 53
rect 1635 -3 2203 53
rect 2259 -3 2827 53
rect 2883 -3 3451 53
rect 3507 -3 4075 53
rect 4131 -3 4699 53
rect 4755 -3 5323 53
rect 5379 -3 5947 53
rect 6003 -3 6571 53
rect 6627 -3 7195 53
rect 7251 -3 7819 53
rect 7875 -3 8443 53
rect 8499 -3 9067 53
rect 9123 -3 9691 53
rect 9747 -3 10315 53
rect 10371 -3 10939 53
rect 10995 -3 11563 53
rect 11619 -3 12187 53
rect 12243 -3 12811 53
rect 12867 -3 13435 53
rect 13491 -3 14059 53
rect 14115 -3 14683 53
rect 14739 -3 15307 53
rect 15363 -3 15931 53
rect 15987 -3 16555 53
rect 16611 -3 17179 53
rect 17235 -3 17803 53
rect 17859 -3 18427 53
rect 18483 -3 19051 53
rect 19107 -3 19675 53
rect 19731 -3 20299 53
rect 20355 -3 20923 53
rect 20979 -3 21547 53
rect 21603 -3 21920 53
rect 33 -8 21920 -3
use subbyte2_precharge_0  subbyte2_precharge_0_0
timestamp 1543373570
transform -1 0 21887 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_1
timestamp 1543373570
transform 1 0 20639 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_2
timestamp 1543373570
transform -1 0 20639 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_3
timestamp 1543373570
transform 1 0 19391 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_4
timestamp 1543373570
transform -1 0 19391 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_5
timestamp 1543373570
transform 1 0 18143 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_6
timestamp 1543373570
transform -1 0 18143 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_7
timestamp 1543373570
transform 1 0 16895 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_8
timestamp 1543373570
transform -1 0 16895 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_9
timestamp 1543373570
transform 1 0 15647 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_10
timestamp 1543373570
transform -1 0 15647 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_11
timestamp 1543373570
transform 1 0 14399 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_12
timestamp 1543373570
transform -1 0 14399 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_13
timestamp 1543373570
transform 1 0 13151 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_14
timestamp 1543373570
transform -1 0 13151 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_15
timestamp 1543373570
transform 1 0 11903 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_16
timestamp 1543373570
transform -1 0 11903 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_17
timestamp 1543373570
transform 1 0 10655 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_18
timestamp 1543373570
transform -1 0 10655 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_19
timestamp 1543373570
transform 1 0 9407 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_20
timestamp 1543373570
transform -1 0 9407 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_21
timestamp 1543373570
transform 1 0 8159 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_22
timestamp 1543373570
transform -1 0 8159 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_23
timestamp 1543373570
transform 1 0 6911 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_24
timestamp 1543373570
transform -1 0 6911 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_25
timestamp 1543373570
transform 1 0 5663 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_26
timestamp 1543373570
transform -1 0 5663 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_27
timestamp 1543373570
transform 1 0 4415 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_28
timestamp 1543373570
transform -1 0 4415 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_29
timestamp 1543373570
transform 1 0 3167 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_30
timestamp 1543373570
transform -1 0 3167 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_31
timestamp 1543373570
transform 1 0 1919 0 1 0
box 0 -8 624 722
use subbyte2_precharge_0  subbyte2_precharge_0_32
timestamp 1543373570
transform -1 0 1919 0 1 0
box 0 -8 624 722
<< labels >>
rlabel metal3 s 33 -8 21920 58 4 en_bar
port 3 nsew
rlabel metal1 s 1825 0 1853 722 4 bl_0
port 5 nsew
rlabel metal1 s 1361 0 1389 722 4 br_0
port 7 nsew
rlabel metal1 s 1985 0 2013 722 4 bl_1
port 9 nsew
rlabel metal1 s 2449 0 2477 722 4 br_1
port 11 nsew
rlabel metal1 s 3073 0 3101 722 4 bl_2
port 13 nsew
rlabel metal1 s 2609 0 2637 722 4 br_2
port 15 nsew
rlabel metal1 s 3233 0 3261 722 4 bl_3
port 17 nsew
rlabel metal1 s 3697 0 3725 722 4 br_3
port 19 nsew
rlabel metal1 s 4321 0 4349 722 4 bl_4
port 21 nsew
rlabel metal1 s 3857 0 3885 722 4 br_4
port 23 nsew
rlabel metal1 s 4481 0 4509 722 4 bl_5
port 25 nsew
rlabel metal1 s 4945 0 4973 722 4 br_5
port 27 nsew
rlabel metal1 s 5569 0 5597 722 4 bl_6
port 29 nsew
rlabel metal1 s 5105 0 5133 722 4 br_6
port 31 nsew
rlabel metal1 s 5729 0 5757 722 4 bl_7
port 33 nsew
rlabel metal1 s 6193 0 6221 722 4 br_7
port 35 nsew
rlabel metal1 s 6817 0 6845 722 4 bl_8
port 37 nsew
rlabel metal1 s 6353 0 6381 722 4 br_8
port 39 nsew
rlabel metal1 s 6977 0 7005 722 4 bl_9
port 41 nsew
rlabel metal1 s 7441 0 7469 722 4 br_9
port 43 nsew
rlabel metal1 s 8065 0 8093 722 4 bl_10
port 45 nsew
rlabel metal1 s 7601 0 7629 722 4 br_10
port 47 nsew
rlabel metal1 s 8225 0 8253 722 4 bl_11
port 49 nsew
rlabel metal1 s 8689 0 8717 722 4 br_11
port 51 nsew
rlabel metal1 s 9313 0 9341 722 4 bl_12
port 53 nsew
rlabel metal1 s 8849 0 8877 722 4 br_12
port 55 nsew
rlabel metal1 s 9473 0 9501 722 4 bl_13
port 57 nsew
rlabel metal1 s 9937 0 9965 722 4 br_13
port 59 nsew
rlabel metal1 s 10561 0 10589 722 4 bl_14
port 61 nsew
rlabel metal1 s 10097 0 10125 722 4 br_14
port 63 nsew
rlabel metal1 s 10721 0 10749 722 4 bl_15
port 65 nsew
rlabel metal1 s 11185 0 11213 722 4 br_15
port 67 nsew
rlabel metal1 s 11809 0 11837 722 4 bl_16
port 69 nsew
rlabel metal1 s 11345 0 11373 722 4 br_16
port 71 nsew
rlabel metal1 s 11969 0 11997 722 4 bl_17
port 73 nsew
rlabel metal1 s 12433 0 12461 722 4 br_17
port 75 nsew
rlabel metal1 s 13057 0 13085 722 4 bl_18
port 77 nsew
rlabel metal1 s 12593 0 12621 722 4 br_18
port 79 nsew
rlabel metal1 s 13217 0 13245 722 4 bl_19
port 81 nsew
rlabel metal1 s 13681 0 13709 722 4 br_19
port 83 nsew
rlabel metal1 s 14305 0 14333 722 4 bl_20
port 85 nsew
rlabel metal1 s 13841 0 13869 722 4 br_20
port 87 nsew
rlabel metal1 s 14465 0 14493 722 4 bl_21
port 89 nsew
rlabel metal1 s 14929 0 14957 722 4 br_21
port 91 nsew
rlabel metal1 s 15553 0 15581 722 4 bl_22
port 93 nsew
rlabel metal1 s 15089 0 15117 722 4 br_22
port 95 nsew
rlabel metal1 s 15713 0 15741 722 4 bl_23
port 97 nsew
rlabel metal1 s 16177 0 16205 722 4 br_23
port 99 nsew
rlabel metal1 s 16801 0 16829 722 4 bl_24
port 101 nsew
rlabel metal1 s 16337 0 16365 722 4 br_24
port 103 nsew
rlabel metal1 s 16961 0 16989 722 4 bl_25
port 105 nsew
rlabel metal1 s 17425 0 17453 722 4 br_25
port 107 nsew
rlabel metal1 s 18049 0 18077 722 4 bl_26
port 109 nsew
rlabel metal1 s 17585 0 17613 722 4 br_26
port 111 nsew
rlabel metal1 s 18209 0 18237 722 4 bl_27
port 113 nsew
rlabel metal1 s 18673 0 18701 722 4 br_27
port 115 nsew
rlabel metal1 s 19297 0 19325 722 4 bl_28
port 117 nsew
rlabel metal1 s 18833 0 18861 722 4 br_28
port 119 nsew
rlabel metal1 s 19457 0 19485 722 4 bl_29
port 121 nsew
rlabel metal1 s 19921 0 19949 722 4 br_29
port 123 nsew
rlabel metal1 s 20545 0 20573 722 4 bl_30
port 125 nsew
rlabel metal1 s 20081 0 20109 722 4 br_30
port 127 nsew
rlabel metal1 s 20705 0 20733 722 4 bl_31
port 129 nsew
rlabel metal1 s 21169 0 21197 722 4 br_31
port 131 nsew
rlabel metal1 s 21793 0 21821 722 4 bl_32
port 133 nsew
rlabel metal1 s 21329 0 21357 722 4 br_32
port 135 nsew
rlabel metal3 s 33 595 21920 661 4 vdd
port 137 nsew
<< properties >>
string FIXED_BBOX 21542 -12 21608 0
<< end >>
