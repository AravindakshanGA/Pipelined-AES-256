
module aes_dec_core (
	clk_clk,
	q_export_readdata,
	reset_reset_n);	

	input		clk_clk;
	output	[63:0]	q_export_readdata;
	input		reset_reset_n;
endmodule
